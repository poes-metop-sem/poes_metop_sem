netcdf poes_nXX_YYYYMMDD_raw {
dimensions:
	time = UNLIMITED ;
variables:
	uint64 time(time) ;
		time:long_name = "milliseconds since 1970-01-01" ;
		time:units = "milliseconds since 1970-01-01" ;
		time:valid_min = 0. ;
		time:_Storage = "chunked" ;
		time:_ChunkSizes = 43200 ;
		time:_DeflateLevel = 9 ;
		time:_Shuffle = "true" ;
		time:_Endianness = "little" ;
	ushort year(time) ;
		year:long_name = "4 digit year" ;
		year:units = "year" ;
		year:valid_range = 1950., 2050. ;
		year:_Storage = "chunked" ;
		year:_ChunkSizes = 43200 ;
		year:_DeflateLevel = 9 ;
		year:_Shuffle = "true" ;
		year:_Endianness = "little" ;
	ushort day(time) ;
		day:long_name = "3 digit day of year" ;
		day:units = "day" ;
		day:valid_range = 0., 366. ;
		day:_Storage = "chunked" ;
		day:_ChunkSizes = 43200 ;
		day:_DeflateLevel = 9 ;
		day:_Shuffle = "true" ;
		day:_Endianness = "little" ;
	uint msec(time) ;
		msec:long_name = "milliseconds of the day" ;
		msec:units = "millisec" ;
		msec:valid_range = 0., 86400000. ;
		msec:_Storage = "chunked" ;
		msec:_ChunkSizes = 43200 ;
		msec:_DeflateLevel = 9 ;
		msec:_Shuffle = "true" ;
		msec:_Endianness = "little" ;
	ubyte satID(time) ;
		satID:long_name = "2 digit number identifying the satellite the data is from" ;
		satID:units = "ID" ;
		satID:valid_range = 0., 20. ;
		satID:_Storage = "chunked" ;
		satID:_ChunkSizes = 43200 ;
		satID:_DeflateLevel = 9 ;
		satID:_Shuffle = "true" ;
	ushort minor_frame(time) ;
		minor_frame:long_name = "minor frame number used to sort data" ;
		minor_frame:units = "frame" ;
		minor_frame:valid_range = 0., 320. ;
		minor_frame:_Storage = "chunked" ;
		minor_frame:_ChunkSizes = 43200 ;
		minor_frame:_DeflateLevel = 9 ;
		minor_frame:_Shuffle = "true" ;
		minor_frame:_Endianness = "little" ;
	ushort major_frame(time) ;
		major_frame:long_name = "major frame number used to sort data" ;
		major_frame:units = "frame" ;
		major_frame:valid_range = 0., 7. ;
		major_frame:_Storage = "chunked" ;
		major_frame:_ChunkSizes = 43200 ;
		major_frame:_DeflateLevel = 9 ;
		major_frame:_Shuffle = "true" ;
		major_frame:_Endianness = "little" ;
	ubyte sat_direction(time) ;
		sat_direction:long_name = "satellite direction 0-North/ 1-South" ;
		sat_direction:units = "" ;
		sat_direction:valid_range = 0., 1. ;
		sat_direction:_Storage = "chunked" ;
		sat_direction:_ChunkSizes = 43200 ;
		sat_direction:_DeflateLevel = 9 ;
		sat_direction:_Shuffle = "true" ;
	float alt(time) ;
		alt:long_name = "altitude of the satellite" ;
		alt:units = "km" ;
		alt:valid_range = 800., 1000. ;
		alt:_Storage = "chunked" ;
		alt:_ChunkSizes = 43200 ;
		alt:_DeflateLevel = 9 ;
		alt:_Shuffle = "true" ;
	float lat(time) ;
		lat:long_name = "latitude of the satellite" ;
		lat:units = "degrees" ;
		lat:valid_range = -90., 90. ;
		lat:_Storage = "chunked" ;
		lat:_ChunkSizes = 43200 ;
		lat:_DeflateLevel = 9 ;
		lat:_Shuffle = "true" ;
	float lon(time) ;
		lon:long_name = "longitude of the satellite" ;
		lon:units = "degrees" ;
		lon:valid_range = 0., 360. ;
		lon:_Storage = "chunked" ;
		lon:_ChunkSizes = 43200 ;
		lon:_DeflateLevel = 9 ;
		lon:_Shuffle = "true" ;
	float mep_pro_tel0_cps_p1(time) ;
		mep_pro_tel0_cps_p1:long_name = "MEPED proton channel 1 ~30-80 keV 0 deg telescope" ;
		mep_pro_tel0_cps_p1:units = "#/s" ;
		mep_pro_tel0_cps_p1:valid_range = 0., 1998848. ;
		mep_pro_tel0_cps_p1:_Storage = "chunked" ;
		mep_pro_tel0_cps_p1:_ChunkSizes = 43200 ;
		mep_pro_tel0_cps_p1:_DeflateLevel = 9 ;
		mep_pro_tel0_cps_p1:_Shuffle = "true" ;
	float mep_pro_tel0_cps_p2(time) ;
		mep_pro_tel0_cps_p2:long_name = "MEPED proton channel 2 ~80-240 keV 0 deg telescope" ;
		mep_pro_tel0_cps_p2:units = "#/s" ;
		mep_pro_tel0_cps_p2:valid_range = 0., 1998848. ;
		mep_pro_tel0_cps_p2:_Storage = "chunked" ;
		mep_pro_tel0_cps_p2:_ChunkSizes = 43200 ;
		mep_pro_tel0_cps_p2:_DeflateLevel = 9 ;
		mep_pro_tel0_cps_p2:_Shuffle = "true" ;
	float mep_pro_tel0_cps_p3(time) ;
		mep_pro_tel0_cps_p3:long_name = "MEPED proton channel 3 ~240-800 keV 0 deg telescope" ;
		mep_pro_tel0_cps_p3:units = "#/s" ;
		mep_pro_tel0_cps_p3:valid_range = 0., 1998848. ;
		mep_pro_tel0_cps_p3:_Storage = "chunked" ;
		mep_pro_tel0_cps_p3:_ChunkSizes = 43200 ;
		mep_pro_tel0_cps_p3:_DeflateLevel = 9 ;
		mep_pro_tel0_cps_p3:_Shuffle = "true" ;
	float mep_pro_tel0_cps_p4(time) ;
		mep_pro_tel0_cps_p4:long_name = "MEPED proton channel 4 ~800-2500 keV 0 deg telescope" ;
		mep_pro_tel0_cps_p4:units = "#/s" ;
		mep_pro_tel0_cps_p4:valid_range = 0., 1998848. ;
		mep_pro_tel0_cps_p4:_Storage = "chunked" ;
		mep_pro_tel0_cps_p4:_ChunkSizes = 43200 ;
		mep_pro_tel0_cps_p4:_DeflateLevel = 9 ;
		mep_pro_tel0_cps_p4:_Shuffle = "true" ;
	float mep_pro_tel0_cps_p5(time) ;
		mep_pro_tel0_cps_p5:long_name = "MEPED proton channel 5 ~2500-6900 keV 0 deg telescope" ;
		mep_pro_tel0_cps_p5:units = "#/s" ;
		mep_pro_tel0_cps_p5:valid_range = 0., 1998848. ;
		mep_pro_tel0_cps_p5:_Storage = "chunked" ;
		mep_pro_tel0_cps_p5:_ChunkSizes = 43200 ;
		mep_pro_tel0_cps_p5:_DeflateLevel = 9 ;
		mep_pro_tel0_cps_p5:_Shuffle = "true" ;
	float mep_pro_tel0_cps_p6(time) ;
		mep_pro_tel0_cps_p6:long_name = "MEPED proton channel 6 ~>6900 keV 0 deg telescope" ;
		mep_pro_tel0_cps_p6:units = "#/s" ;
		mep_pro_tel0_cps_p6:valid_range = 0., 1998848. ;
		mep_pro_tel0_cps_p6:_Storage = "chunked" ;
		mep_pro_tel0_cps_p6:_ChunkSizes = 43200 ;
		mep_pro_tel0_cps_p6:_DeflateLevel = 9 ;
		mep_pro_tel0_cps_p6:_Shuffle = "true" ;
	float mep_pro_tel90_cps_p1(time) ;
		mep_pro_tel90_cps_p1:long_name = "MEPED proton channel 1 ~30-80 keV 90 deg telescope" ;
		mep_pro_tel90_cps_p1:units = "#/s" ;
		mep_pro_tel90_cps_p1:valid_range = 0., 1998848. ;
		mep_pro_tel90_cps_p1:_Storage = "chunked" ;
		mep_pro_tel90_cps_p1:_ChunkSizes = 43200 ;
		mep_pro_tel90_cps_p1:_DeflateLevel = 9 ;
		mep_pro_tel90_cps_p1:_Shuffle = "true" ;
	float mep_pro_tel90_cps_p2(time) ;
		mep_pro_tel90_cps_p2:long_name = "MEPED proton channel 2 ~80-240 keV 90 deg telescope" ;
		mep_pro_tel90_cps_p2:units = "#/s" ;
		mep_pro_tel90_cps_p2:valid_range = 0., 1998848. ;
		mep_pro_tel90_cps_p2:_Storage = "chunked" ;
		mep_pro_tel90_cps_p2:_ChunkSizes = 43200 ;
		mep_pro_tel90_cps_p2:_DeflateLevel = 9 ;
		mep_pro_tel90_cps_p2:_Shuffle = "true" ;
	float mep_pro_tel90_cps_p3(time) ;
		mep_pro_tel90_cps_p3:long_name = "MEPED proton channel 3 ~240-800 keV 90 deg telescope" ;
		mep_pro_tel90_cps_p3:units = "#/s" ;
		mep_pro_tel90_cps_p3:valid_range = 0., 1998848. ;
		mep_pro_tel90_cps_p3:_Storage = "chunked" ;
		mep_pro_tel90_cps_p3:_ChunkSizes = 43200 ;
		mep_pro_tel90_cps_p3:_DeflateLevel = 9 ;
		mep_pro_tel90_cps_p3:_Shuffle = "true" ;
	float mep_pro_tel90_cps_p4(time) ;
		mep_pro_tel90_cps_p4:long_name = "MEPED proton channel 4 ~800-2500 keV 90 deg telescope" ;
		mep_pro_tel90_cps_p4:units = "#/s" ;
		mep_pro_tel90_cps_p4:valid_range = 0., 1998848. ;
		mep_pro_tel90_cps_p4:_Storage = "chunked" ;
		mep_pro_tel90_cps_p4:_ChunkSizes = 43200 ;
		mep_pro_tel90_cps_p4:_DeflateLevel = 9 ;
		mep_pro_tel90_cps_p4:_Shuffle = "true" ;
	float mep_pro_tel90_cps_p5(time) ;
		mep_pro_tel90_cps_p5:long_name = "MEPED proton channel 5 ~2500-6900 keV 90 deg telescope" ;
		mep_pro_tel90_cps_p5:units = "#/s" ;
		mep_pro_tel90_cps_p5:valid_range = 0., 1998848. ;
		mep_pro_tel90_cps_p5:_Storage = "chunked" ;
		mep_pro_tel90_cps_p5:_ChunkSizes = 43200 ;
		mep_pro_tel90_cps_p5:_DeflateLevel = 9 ;
		mep_pro_tel90_cps_p5:_Shuffle = "true" ;
	float mep_pro_tel90_cps_p6(time) ;
		mep_pro_tel90_cps_p6:long_name = "MEPED proton channel 6 ~>6900 keV 90 degree telescope" ;
		mep_pro_tel90_cps_p6:units = "#/s" ;
		mep_pro_tel90_cps_p6:valid_range = 0., 1998848. ;
		mep_pro_tel90_cps_p6:_Storage = "chunked" ;
		mep_pro_tel90_cps_p6:_ChunkSizes = 43200 ;
		mep_pro_tel90_cps_p6:_DeflateLevel = 9 ;
		mep_pro_tel90_cps_p6:_Shuffle = "true" ;
	float mep_ele_tel0_cps_e1(time) ;
		mep_ele_tel0_cps_e1:long_name = "MEPED electron channel 1 ~>30 keV #/s 0 deg telescope" ;
		mep_ele_tel0_cps_e1:units = "#/s" ;
		mep_ele_tel0_cps_e1:valid_range = 0., 1998848. ;
		mep_ele_tel0_cps_e1:_Storage = "chunked" ;
		mep_ele_tel0_cps_e1:_ChunkSizes = 43200 ;
		mep_ele_tel0_cps_e1:_DeflateLevel = 9 ;
		mep_ele_tel0_cps_e1:_Shuffle = "true" ;
	float mep_ele_tel0_cps_e2(time) ;
		mep_ele_tel0_cps_e2:long_name = "MEPED electron channel 2 ~>100 keV #/s 0 deg telescope" ;
		mep_ele_tel0_cps_e2:units = "#/s" ;
		mep_ele_tel0_cps_e2:valid_range = 0., 1998848. ;
		mep_ele_tel0_cps_e2:_Storage = "chunked" ;
		mep_ele_tel0_cps_e2:_ChunkSizes = 43200 ;
		mep_ele_tel0_cps_e2:_DeflateLevel = 9 ;
		mep_ele_tel0_cps_e2:_Shuffle = "true" ;
	float mep_ele_tel0_cps_e3(time) ;
		mep_ele_tel0_cps_e3:long_name = "MEPED electron channel 3 ~>300 keV #/s 0 deg telescope" ;
		mep_ele_tel0_cps_e3:units = "#/s" ;
		mep_ele_tel0_cps_e3:valid_range = 0., 1998848. ;
		mep_ele_tel0_cps_e3:_Storage = "chunked" ;
		mep_ele_tel0_cps_e3:_ChunkSizes = 43200 ;
		mep_ele_tel0_cps_e3:_DeflateLevel = 9 ;
		mep_ele_tel0_cps_e3:_Shuffle = "true" ;
	float mep_ele_tel90_cps_e1(time) ;
		mep_ele_tel90_cps_e1:long_name = "MEPED electron channel 1 ~>30 keV #/s 90 deg telescope" ;
		mep_ele_tel90_cps_e1:units = "#/s" ;
		mep_ele_tel90_cps_e1:valid_range = 0., 1998848. ;
		mep_ele_tel90_cps_e1:_Storage = "chunked" ;
		mep_ele_tel90_cps_e1:_ChunkSizes = 43200 ;
		mep_ele_tel90_cps_e1:_DeflateLevel = 9 ;
		mep_ele_tel90_cps_e1:_Shuffle = "true" ;
	float mep_ele_tel90_cps_e2(time) ;
		mep_ele_tel90_cps_e2:long_name = "MEPED electron channel 2 ~>100 keV #/s 90 deg telescope" ;
		mep_ele_tel90_cps_e2:units = "#/s" ;
		mep_ele_tel90_cps_e2:valid_range = 0., 1998848. ;
		mep_ele_tel90_cps_e2:_Storage = "chunked" ;
		mep_ele_tel90_cps_e2:_ChunkSizes = 43200 ;
		mep_ele_tel90_cps_e2:_DeflateLevel = 9 ;
		mep_ele_tel90_cps_e2:_Shuffle = "true" ;
	float mep_ele_tel90_cps_e3(time) ;
		mep_ele_tel90_cps_e3:long_name = "MEPED electron channel 3 ~>300 keV #/s 90 deg telescope" ;
		mep_ele_tel90_cps_e3:units = "#/s" ;
		mep_ele_tel90_cps_e3:valid_range = 0., 1998848. ;
		mep_ele_tel90_cps_e3:_Storage = "chunked" ;
		mep_ele_tel90_cps_e3:_ChunkSizes = 43200 ;
		mep_ele_tel90_cps_e3:_DeflateLevel = 9 ;
		mep_ele_tel90_cps_e3:_Shuffle = "true" ;
	float mep_omni_cps_p6(time) ;
		mep_omni_cps_p6:long_name = "MEPED proton channel p6 ~>16 MeV omnidirectional telescope" ;
		mep_omni_cps_p6:units = "#/s" ;
		mep_omni_cps_p6:valid_range = 0., 1998848. ;
		mep_omni_cps_p6:_Storage = "chunked" ;
		mep_omni_cps_p6:_ChunkSizes = 43200 ;
		mep_omni_cps_p6:_DeflateLevel = 9 ;
		mep_omni_cps_p6:_Shuffle = "true" ;
	float mep_omni_cps_p7(time) ;
		mep_omni_cps_p7:long_name = "MEPED proton channel p7 ~>35 MeV omnidirectional telescope" ;
		mep_omni_cps_p7:units = "#/s" ;
		mep_omni_cps_p7:valid_range = 0., 1998848. ;
		mep_omni_cps_p7:_Storage = "chunked" ;
		mep_omni_cps_p7:_ChunkSizes = 43200 ;
		mep_omni_cps_p7:_DeflateLevel = 9 ;
		mep_omni_cps_p7:_Shuffle = "true" ;
	float mep_omni_cps_p8(time) ;
		mep_omni_cps_p8:long_name = "MEPED proton channel p8 ~>70 MeV omnidirectional telescope" ;
		mep_omni_cps_p8:units = "#/s" ;
		mep_omni_cps_p8:valid_range = 0., 1998848. ;
		mep_omni_cps_p8:_Storage = "chunked" ;
		mep_omni_cps_p8:_ChunkSizes = 43200 ;
		mep_omni_cps_p8:_DeflateLevel = 9 ;
		mep_omni_cps_p8:_Shuffle = "true" ;
	float mep_omni_cps_p9(time) ;
		mep_omni_cps_p9:long_name = "MEPED proton channel p9 ~>140 MeV omnidirectional telescope" ;
		mep_omni_cps_p9:units = "#/s" ;
		mep_omni_cps_p9:valid_range = 0., 1998848. ;
		mep_omni_cps_p9:_Storage = "chunked" ;
		mep_omni_cps_p9:_ChunkSizes = 43200 ;
		mep_omni_cps_p9:_DeflateLevel = 9 ;
		mep_omni_cps_p9:_Shuffle = "true" ;
	float ted_ele_tel0_cps_4(time) ;
		ted_ele_tel0_cps_4:long_name = "TED electron energy band 4 0 deg telescope" ;
		ted_ele_tel0_cps_4:units = "counts" ;
		ted_ele_tel0_cps_4:valid_range = 0., 1998848. ;
		ted_ele_tel0_cps_4:_Storage = "chunked" ;
		ted_ele_tel0_cps_4:_ChunkSizes = 43200 ;
		ted_ele_tel0_cps_4:_DeflateLevel = 9 ;
		ted_ele_tel0_cps_4:_Shuffle = "true" ;
	float ted_ele_tel0_cps_8(time) ;
		ted_ele_tel0_cps_8:long_name = "TED electron energy band 8 0 deg telescope" ;
		ted_ele_tel0_cps_8:units = "counts" ;
		ted_ele_tel0_cps_8:valid_range = 0., 1998848. ;
		ted_ele_tel0_cps_8:_Storage = "chunked" ;
		ted_ele_tel0_cps_8:_ChunkSizes = 43200 ;
		ted_ele_tel0_cps_8:_DeflateLevel = 9 ;
		ted_ele_tel0_cps_8:_Shuffle = "true" ;
	float ted_ele_tel0_cps_11(time) ;
		ted_ele_tel0_cps_11:long_name = "TED electron energy band 11 0 deg telescope" ;
		ted_ele_tel0_cps_11:units = "counts" ;
		ted_ele_tel0_cps_11:valid_range = 0., 1998848. ;
		ted_ele_tel0_cps_11:_Storage = "chunked" ;
		ted_ele_tel0_cps_11:_ChunkSizes = 43200 ;
		ted_ele_tel0_cps_11:_DeflateLevel = 9 ;
		ted_ele_tel0_cps_11:_Shuffle = "true" ;
	float ted_ele_tel0_cps_14(time) ;
		ted_ele_tel0_cps_14:long_name = "TED electron energy band 14 0 deg telescope" ;
		ted_ele_tel0_cps_14:units = "counts" ;
		ted_ele_tel0_cps_14:valid_range = 0., 1998848. ;
		ted_ele_tel0_cps_14:_Storage = "chunked" ;
		ted_ele_tel0_cps_14:_ChunkSizes = 43200 ;
		ted_ele_tel0_cps_14:_DeflateLevel = 9 ;
		ted_ele_tel0_cps_14:_Shuffle = "true" ;
	float ted_ele_tel30_cps_4(time) ;
		ted_ele_tel30_cps_4:long_name = "TED electron energy band 4 30 deg telescope" ;
		ted_ele_tel30_cps_4:units = "counts" ;
		ted_ele_tel30_cps_4:valid_range = 0., 1998848. ;
		ted_ele_tel30_cps_4:_Storage = "chunked" ;
		ted_ele_tel30_cps_4:_ChunkSizes = 43200 ;
		ted_ele_tel30_cps_4:_DeflateLevel = 9 ;
		ted_ele_tel30_cps_4:_Shuffle = "true" ;
	float ted_ele_tel30_cps_8(time) ;
		ted_ele_tel30_cps_8:long_name = "TED electron energy band 8 30 deg telescope" ;
		ted_ele_tel30_cps_8:units = "counts" ;
		ted_ele_tel30_cps_8:valid_range = 0., 1998848. ;
		ted_ele_tel30_cps_8:_Storage = "chunked" ;
		ted_ele_tel30_cps_8:_ChunkSizes = 43200 ;
		ted_ele_tel30_cps_8:_DeflateLevel = 9 ;
		ted_ele_tel30_cps_8:_Shuffle = "true" ;
	float ted_ele_tel30_cps_11(time) ;
		ted_ele_tel30_cps_11:long_name = "TED electron energy band 11 30 deg telescope" ;
		ted_ele_tel30_cps_11:units = "counts" ;
		ted_ele_tel30_cps_11:valid_range = 0., 1998848. ;
		ted_ele_tel30_cps_11:_Storage = "chunked" ;
		ted_ele_tel30_cps_11:_ChunkSizes = 43200 ;
		ted_ele_tel30_cps_11:_DeflateLevel = 9 ;
		ted_ele_tel30_cps_11:_Shuffle = "true" ;
	float ted_ele_tel30_cps_14(time) ;
		ted_ele_tel30_cps_14:long_name = "TED electron energy band 14 30 deg telescope" ;
		ted_ele_tel30_cps_14:units = "counts" ;
		ted_ele_tel30_cps_14:valid_range = 0., 1998848. ;
		ted_ele_tel30_cps_14:_Storage = "chunked" ;
		ted_ele_tel30_cps_14:_ChunkSizes = 43200 ;
		ted_ele_tel30_cps_14:_DeflateLevel = 9 ;
		ted_ele_tel30_cps_14:_Shuffle = "true" ;
	float ted_pro_tel0_cps_4(time) ;
		ted_pro_tel0_cps_4:long_name = "TED proton energy band 4 0 deg telescope" ;
		ted_pro_tel0_cps_4:units = "counts" ;
		ted_pro_tel0_cps_4:valid_range = 0., 1998848. ;
		ted_pro_tel0_cps_4:_Storage = "chunked" ;
		ted_pro_tel0_cps_4:_ChunkSizes = 43200 ;
		ted_pro_tel0_cps_4:_DeflateLevel = 9 ;
		ted_pro_tel0_cps_4:_Shuffle = "true" ;
	float ted_pro_tel0_cps_8(time) ;
		ted_pro_tel0_cps_8:long_name = "TED proton energy band 8 0 deg telescope" ;
		ted_pro_tel0_cps_8:units = "counts" ;
		ted_pro_tel0_cps_8:valid_range = 0., 1998848. ;
		ted_pro_tel0_cps_8:_Storage = "chunked" ;
		ted_pro_tel0_cps_8:_ChunkSizes = 43200 ;
		ted_pro_tel0_cps_8:_DeflateLevel = 9 ;
		ted_pro_tel0_cps_8:_Shuffle = "true" ;
	float ted_pro_tel0_cps_11(time) ;
		ted_pro_tel0_cps_11:long_name = "TED proton energy band 11 0 deg telescope" ;
		ted_pro_tel0_cps_11:units = "counts" ;
		ted_pro_tel0_cps_11:valid_range = 0., 1998848. ;
		ted_pro_tel0_cps_11:_Storage = "chunked" ;
		ted_pro_tel0_cps_11:_ChunkSizes = 43200 ;
		ted_pro_tel0_cps_11:_DeflateLevel = 9 ;
		ted_pro_tel0_cps_11:_Shuffle = "true" ;
	float ted_pro_tel0_cps_14(time) ;
		ted_pro_tel0_cps_14:long_name = "TED proton energy band 14 0 deg telescope" ;
		ted_pro_tel0_cps_14:units = "counts" ;
		ted_pro_tel0_cps_14:valid_range = 0., 1998848. ;
		ted_pro_tel0_cps_14:_Storage = "chunked" ;
		ted_pro_tel0_cps_14:_ChunkSizes = 43200 ;
		ted_pro_tel0_cps_14:_DeflateLevel = 9 ;
		ted_pro_tel0_cps_14:_Shuffle = "true" ;
	float ted_pro_tel30_cps_4(time) ;
		ted_pro_tel30_cps_4:long_name = "TED proton energy band 4 30 deg telescope" ;
		ted_pro_tel30_cps_4:units = "counts" ;
		ted_pro_tel30_cps_4:valid_range = 0., 1998848. ;
		ted_pro_tel30_cps_4:_Storage = "chunked" ;
		ted_pro_tel30_cps_4:_ChunkSizes = 43200 ;
		ted_pro_tel30_cps_4:_DeflateLevel = 9 ;
		ted_pro_tel30_cps_4:_Shuffle = "true" ;
	float ted_pro_tel30_cps_8(time) ;
		ted_pro_tel30_cps_8:long_name = "TED proton energy band 8 30 deg telescope" ;
		ted_pro_tel30_cps_8:units = "counts" ;
		ted_pro_tel30_cps_8:valid_range = 0., 1998848. ;
		ted_pro_tel30_cps_8:_Storage = "chunked" ;
		ted_pro_tel30_cps_8:_ChunkSizes = 43200 ;
		ted_pro_tel30_cps_8:_DeflateLevel = 9 ;
		ted_pro_tel30_cps_8:_Shuffle = "true" ;
	float ted_pro_tel30_cps_11(time) ;
		ted_pro_tel30_cps_11:long_name = "TED proton energy band 11 30 deg telescope" ;
		ted_pro_tel30_cps_11:units = "counts" ;
		ted_pro_tel30_cps_11:valid_range = 0., 1998848. ;
		ted_pro_tel30_cps_11:_Storage = "chunked" ;
		ted_pro_tel30_cps_11:_ChunkSizes = 43200 ;
		ted_pro_tel30_cps_11:_DeflateLevel = 9 ;
		ted_pro_tel30_cps_11:_Shuffle = "true" ;
	float ted_pro_tel30_cps_14(time) ;
		ted_pro_tel30_cps_14:long_name = "TED proton energy band 14 30 deg telescope" ;
		ted_pro_tel30_cps_14:units = "counts" ;
		ted_pro_tel30_cps_14:valid_range = 0., 1998848. ;
		ted_pro_tel30_cps_14:_Storage = "chunked" ;
		ted_pro_tel30_cps_14:_ChunkSizes = 43200 ;
		ted_pro_tel30_cps_14:_DeflateLevel = 9 ;
		ted_pro_tel30_cps_14:_Shuffle = "true" ;
	float ted_ele_tel0_low_eflux_cps(time) ;
		ted_ele_tel0_low_eflux_cps:long_name = "TED electron (50eV-1 keV) 0 deg telescope energy flux" ;
		ted_ele_tel0_low_eflux_cps:units = "counts" ;
		ted_ele_tel0_low_eflux_cps:valid_range = 0., 1998848. ;
		ted_ele_tel0_low_eflux_cps:_Storage = "chunked" ;
		ted_ele_tel0_low_eflux_cps:_ChunkSizes = 43200 ;
		ted_ele_tel0_low_eflux_cps:_DeflateLevel = 9 ;
		ted_ele_tel0_low_eflux_cps:_Shuffle = "true" ;
	float ted_ele_tel30_low_eflux_cps(time) ;
		ted_ele_tel30_low_eflux_cps:long_name = "TED electron (50eV-1 keV) 30 deg telescope energy flux" ;
		ted_ele_tel30_low_eflux_cps:units = "counts" ;
		ted_ele_tel30_low_eflux_cps:valid_range = 0., 1998848. ;
		ted_ele_tel30_low_eflux_cps:_Storage = "chunked" ;
		ted_ele_tel30_low_eflux_cps:_ChunkSizes = 43200 ;
		ted_ele_tel30_low_eflux_cps:_DeflateLevel = 9 ;
		ted_ele_tel30_low_eflux_cps:_Shuffle = "true" ;
	float ted_ele_tel0_hi_eflux_cps(time) ;
		ted_ele_tel0_hi_eflux_cps:long_name = "TED electron (1-20 keV) 0 deg telescope energy flux" ;
		ted_ele_tel0_hi_eflux_cps:units = "counts" ;
		ted_ele_tel0_hi_eflux_cps:valid_range = 0., 1998848. ;
		ted_ele_tel0_hi_eflux_cps:_Storage = "chunked" ;
		ted_ele_tel0_hi_eflux_cps:_ChunkSizes = 43200 ;
		ted_ele_tel0_hi_eflux_cps:_DeflateLevel = 9 ;
		ted_ele_tel0_hi_eflux_cps:_Shuffle = "true" ;
	float ted_ele_tel30_hi_eflux_cps(time) ;
		ted_ele_tel30_hi_eflux_cps:long_name = "TED electron (1-20 keV)  30 deg telescope energy flux" ;
		ted_ele_tel30_hi_eflux_cps:units = "counts" ;
		ted_ele_tel30_hi_eflux_cps:valid_range = 0., 1998848. ;
		ted_ele_tel30_hi_eflux_cps:_Storage = "chunked" ;
		ted_ele_tel30_hi_eflux_cps:_ChunkSizes = 43200 ;
		ted_ele_tel30_hi_eflux_cps:_DeflateLevel = 9 ;
		ted_ele_tel30_hi_eflux_cps:_Shuffle = "true" ;
	float ted_pro_tel0_low_eflux_cps(time) ;
		ted_pro_tel0_low_eflux_cps:long_name = "TED proton (50eV-1 keV) 0 deg telescope energy flux" ;
		ted_pro_tel0_low_eflux_cps:units = "counts" ;
		ted_pro_tel0_low_eflux_cps:valid_range = 0., 1998848. ;
		ted_pro_tel0_low_eflux_cps:_Storage = "chunked" ;
		ted_pro_tel0_low_eflux_cps:_ChunkSizes = 43200 ;
		ted_pro_tel0_low_eflux_cps:_DeflateLevel = 9 ;
		ted_pro_tel0_low_eflux_cps:_Shuffle = "true" ;
	float ted_pro_tel30_low_eflux_cps(time) ;
		ted_pro_tel30_low_eflux_cps:long_name = "TEDproton (50eV-1 keV) 30 deg telescope energy flux" ;
		ted_pro_tel30_low_eflux_cps:units = "counts" ;
		ted_pro_tel30_low_eflux_cps:valid_range = 0., 1998848. ;
		ted_pro_tel30_low_eflux_cps:_Storage = "chunked" ;
		ted_pro_tel30_low_eflux_cps:_ChunkSizes = 43200 ;
		ted_pro_tel30_low_eflux_cps:_DeflateLevel = 9 ;
		ted_pro_tel30_low_eflux_cps:_Shuffle = "true" ;
	float ted_pro_tel0_hi_eflux_cps(time) ;
		ted_pro_tel0_hi_eflux_cps:long_name = "TED proton (1-20 keV)  0 deg telescope energy flux" ;
		ted_pro_tel0_hi_eflux_cps:units = "counts" ;
		ted_pro_tel0_hi_eflux_cps:valid_range = 0., 1998848. ;
		ted_pro_tel0_hi_eflux_cps:_Storage = "chunked" ;
		ted_pro_tel0_hi_eflux_cps:_ChunkSizes = 43200 ;
		ted_pro_tel0_hi_eflux_cps:_DeflateLevel = 9 ;
		ted_pro_tel0_hi_eflux_cps:_Shuffle = "true" ;
	float ted_pro_tel30_hi_eflux_cps(time) ;
		ted_pro_tel30_hi_eflux_cps:long_name = "TED proton (1-20 keV)  30 deg telescope energy flux" ;
		ted_pro_tel30_hi_eflux_cps:units = "counts" ;
		ted_pro_tel30_hi_eflux_cps:valid_range = 0., 1998848. ;
		ted_pro_tel30_hi_eflux_cps:_Storage = "chunked" ;
		ted_pro_tel30_hi_eflux_cps:_ChunkSizes = 43200 ;
		ted_pro_tel30_hi_eflux_cps:_DeflateLevel = 9 ;
		ted_pro_tel30_hi_eflux_cps:_Shuffle = "true" ;
	float microA_V(time) ;
		microA_V:long_name = "microprocessor A Voltage [+5 V nominal]" ;
		microA_V:units = "V" ;
		microA_V:_Storage = "chunked" ;
		microA_V:_ChunkSizes = 43200 ;
		microA_V:_DeflateLevel = 9 ;
		microA_V:_Shuffle = "true" ;
	float microB_V(time) ;
		microB_V:long_name = "microprocessor B Voltage [+5 V nominal]" ;
		microB_V:units = "V" ;
		microB_V:_Storage = "chunked" ;
		microB_V:_ChunkSizes = 43200 ;
		microB_V:_DeflateLevel = 9 ;
		microB_V:_Shuffle = "true" ;
	float DPU_V(time) ;
		DPU_V:long_name = "DPU voltage [+5 V nominal]" ;
		DPU_V:units = "V" ;
		DPU_V:_Storage = "chunked" ;
		DPU_V:_ChunkSizes = 43200 ;
		DPU_V:_DeflateLevel = 9 ;
		DPU_V:_Shuffle = "true" ;
	float MEPED_V(time) ;
		MEPED_V:long_name = "MEPED voltage [+5 V nominal]" ;
		MEPED_V:units = "V" ;
		MEPED_V:_Storage = "chunked" ;
		MEPED_V:_ChunkSizes = 43200 ;
		MEPED_V:_DeflateLevel = 9 ;
		MEPED_V:_Shuffle = "true" ;
	float ted_V(time) ;
		ted_V:long_name = "TED voltage [+5 V nominal]" ;
		ted_V:units = "V" ;
		ted_V:_Storage = "chunked" ;
		ted_V:_ChunkSizes = 43200 ;
		ted_V:_DeflateLevel = 9 ;
		ted_V:_Shuffle = "true" ;
	float ted_sweepV(time) ;
		ted_sweepV:long_name = "TED sweep voltage" ;
		ted_sweepV:units = "V" ;
		ted_sweepV:_Storage = "chunked" ;
		ted_sweepV:_ChunkSizes = 43200 ;
		ted_sweepV:_DeflateLevel = 9 ;
		ted_sweepV:_Shuffle = "true" ;
	float ted_electron_CEM_V(time) ;
		ted_electron_CEM_V:long_name = "TED electron CEM voltage" ;
		ted_electron_CEM_V:units = "V" ;
		ted_electron_CEM_V:_Storage = "chunked" ;
		ted_electron_CEM_V:_ChunkSizes = 43200 ;
		ted_electron_CEM_V:_DeflateLevel = 9 ;
		ted_electron_CEM_V:_Shuffle = "true" ;
	float ted_proton_CEM_V(time) ;
		ted_proton_CEM_V:long_name = "TED proton CEM voltage" ;
		ted_proton_CEM_V:units = "V" ;
		ted_proton_CEM_V:_Storage = "chunked" ;
		ted_proton_CEM_V:_ChunkSizes = 43200 ;
		ted_proton_CEM_V:_DeflateLevel = 9 ;
		ted_proton_CEM_V:_Shuffle = "true" ;
	float mep_omni_biase_V(time) ;
		mep_omni_biase_V:long_name = "MEPED omni bias voltage" ;
		mep_omni_biase_V:units = "V" ;
		mep_omni_biase_V:_Storage = "chunked" ;
		mep_omni_biase_V:_ChunkSizes = 43200 ;
		mep_omni_biase_V:_DeflateLevel = 9 ;
		mep_omni_biase_V:_Shuffle = "true" ;
	float mep_circuit_temp(time) ;
		mep_circuit_temp:long_name = "MEPED electronic circuit temperature" ;
		mep_circuit_temp:units = "K" ;
		mep_circuit_temp:_Storage = "chunked" ;
		mep_circuit_temp:_ChunkSizes = 43200 ;
		mep_circuit_temp:_DeflateLevel = 9 ;
		mep_circuit_temp:_Shuffle = "true" ;
	float mep_proton_tel_temp(time) ;
		mep_proton_tel_temp:long_name = "MEPED proton telescope temperature" ;
		mep_proton_tel_temp:units = "K" ;
		mep_proton_tel_temp:_Storage = "chunked" ;
		mep_proton_tel_temp:_ChunkSizes = 43200 ;
		mep_proton_tel_temp:_DeflateLevel = 9 ;
		mep_proton_tel_temp:_Shuffle = "true" ;
	float TED_temp(time) ;
		TED_temp:long_name = "TED temperature" ;
		TED_temp:units = "K" ;
		TED_temp:_Storage = "chunked" ;
		TED_temp:_ChunkSizes = 43200 ;
		TED_temp:_DeflateLevel = 9 ;
		TED_temp:_Shuffle = "true" ;
	float DPU_temp(time) ;
		DPU_temp:long_name = "DPU temperature" ;
		DPU_temp:units = "K" ;
		DPU_temp:_Storage = "chunked" ;
		DPU_temp:_ChunkSizes = 43200 ;
		DPU_temp:_DeflateLevel = 9 ;
		DPU_temp:_Shuffle = "true" ;
	float HK_data(time) ;
		HK_data:long_name = "housekeeping data" ;
		HK_data:units = "variable" ;
		HK_data:_Storage = "chunked" ;
		HK_data:_ChunkSizes = 43200 ;
		HK_data:_DeflateLevel = 9 ;
		HK_data:_Shuffle = "true" ;
	byte HK_key(time) ;
		HK_key:long_name = "key for interpreting housekeeping data" ;
		HK_key:units = "key value" ;
		HK_key:_Storage = "chunked" ;
		HK_key:_ChunkSizes = 43200 ;
		HK_key:_DeflateLevel = 9 ;
		HK_key:_Shuffle = "true" ;
	byte ted_ele_PHD_level(time) ;
		ted_ele_PHD_level:long_name = "TED electron pulse height discriminator level" ;
		ted_ele_PHD_level:units = "level" ;
		ted_ele_PHD_level:valid_range = 0., 3. ;
		ted_ele_PHD_level:_Storage = "chunked" ;
		ted_ele_PHD_level:_ChunkSizes = 43200 ;
		ted_ele_PHD_level:_DeflateLevel = 9 ;
		ted_ele_PHD_level:_Shuffle = "true" ;
	byte ted_pro_PHD_level(time) ;
		ted_pro_PHD_level:long_name = "TED proton pulse height discriminator level" ;
		ted_pro_PHD_level:units = "level" ;
		ted_pro_PHD_level:valid_range = 0., 3. ;
		ted_pro_PHD_level:_Storage = "chunked" ;
		ted_pro_PHD_level:_ChunkSizes = 43200 ;
		ted_pro_PHD_level:_DeflateLevel = 9 ;
		ted_pro_PHD_level:_Shuffle = "true" ;
	byte ted_IFC_on(time) ;
		ted_IFC_on:long_name = "TED IFC flag (0 off 1 on)" ;
		ted_IFC_on:units = "on/off" ;
		ted_IFC_on:valid_range = 0., 1. ;
		ted_IFC_on:_Storage = "chunked" ;
		ted_IFC_on:_ChunkSizes = 43200 ;
		ted_IFC_on:_DeflateLevel = 9 ;
		ted_IFC_on:_Shuffle = "true" ;
                ted_IFC_on:_FillValue = -1 ;
	byte mep_IFC_on(time) ;
		mep_IFC_on:long_name = "MEPED IFC flag (0 off 1 on)" ;
		mep_IFC_on:units = "on/off" ;
		mep_IFC_on:valid_range = 0., 1. ;
		mep_IFC_on:_Storage = "chunked" ;
		mep_IFC_on:_ChunkSizes = 43200 ;
		mep_IFC_on:_DeflateLevel = 9 ;
		mep_IFC_on:_Shuffle = "true" ;
                mep_IFC_on:_FillValue = -1 ;
	byte ted_ele_HV_step(time) ;
		ted_ele_HV_step:long_name = "TED electron high voltage step" ;
		ted_ele_HV_step:units = "step" ;
		ted_ele_HV_step:valid_range = 0., 7. ;
		ted_ele_HV_step:_Storage = "chunked" ;
		ted_ele_HV_step:_ChunkSizes = 43200 ;
		ted_ele_HV_step:_DeflateLevel = 9 ;
		ted_ele_HV_step:_Shuffle = "true" ;
	byte ted_pro_HV_step(time) ;
		ted_pro_HV_step:long_name = "TED proton high voltage step" ;
		ted_pro_HV_step:units = "step" ;
		ted_pro_HV_step:valid_range = 0., 7. ;
		ted_pro_HV_step:_Storage = "chunked" ;
		ted_pro_HV_step:_ChunkSizes = 43200 ;
		ted_pro_HV_step:_DeflateLevel = 9 ;
		ted_pro_HV_step:_Shuffle = "true" ;

// global attributes:
		:title = "POES/MetOp: Particle Precipitation (These data have known contamination problems. Please consult provider for usage recommendations.)" ;
		:naming_authority = "" ;
		:time_coverage_duration = "1day" ;
		:time_coverage_resolution = "2sec" ;
		:geospatial_lat_min = "-90" ;
		:geospatial_lat_max = "90" ;
		:geospatial_lat_unit = "degrees" ;
		:geospatial_lon_min = "0" ;
		:geospatial_lon_max = "360" ;
		:geospatial_lon_units = "degrees East" ;
		:geospatial_vertical_min = "850" ;
		:geospatial_vertical_max = "850" ;
		:geospatial_vertical_units = "km" ;
		:geospatial_vertical_positive = "up" ;
		:point_of_contact = "" ;
		:institution = "" ;
		:creator = "" ;
		:creator_url = "" ;
		:creator_email = "" ;
		:publisher_name = "" ;
		:publisher_url = "" ;
		:publisher_email = "" ;
		:release = "Public Release" ;
		:description = "POES/MetOp SEM-2 Data" ;
		:summary = "The POES/MetOp SEM-2 data provide information about the particle radiation surrounding Earth and its effects on the atmosphere" ;
		:keywords_vocabulary = "Earth Science > Sun-earth Interactions > Ionosphere/Magnetosphere Particles > Electron Flux,Earth Science > Sun-earth Interactions > Ionosphere/Magnetosphere Particles " ;
		:comment = "Every effort has been made to provide the highest quality data but the instruments have known inherent limitations. Please contact the data provider for information on how to properly use the data." ;
		:license = "Public" ;
		:Project = "POES/MetOp" ;
		:processing_level = "Level 2, calibrated fluxes" ;
		:_Format = "netCDF-4" ;
}
