netcdf poes_nXX_YYYYMMDD_proc {
dimensions:
	time = UNLIMITED ;
variables:
	uint64 time(time) ;
		time:long_name = "milliseconds since 1970-01-01" ;
		time:units = "milliseconds since 1970-01-01" ;
		time:valid_min = 0. ;
		time:_Storage = "chunked" ;
		time:_ChunkSizes = 43200 ;
		time:_DeflateLevel = 9 ;
		time:_Shuffle = "true" ;
		time:_Endianness = "little" ;
	ushort year(time) ;
		year:long_name = "4 digit year" ;
		year:units = "year" ;
		year:valid_range = 1950., 2050. ;
		year:_Storage = "chunked" ;
		year:_ChunkSizes = 43200 ;
		year:_DeflateLevel = 9 ;
		year:_Shuffle = "true" ;
		year:_Endianness = "little" ;
	ushort day(time) ;
		day:long_name = "3 digit day of year" ;
		day:units = "day" ;
		day:valid_range = 0., 366. ;
		day:_Storage = "chunked" ;
		day:_ChunkSizes = 43200 ;
		day:_DeflateLevel = 9 ;
		day:_Shuffle = "true" ;
		day:_Endianness = "little" ;
	uint msec(time) ;
		msec:long_name = "milliseconds of the day" ;
		msec:units = "millisec" ;
		msec:valid_range = 0., 86400000. ;
		msec:_Storage = "chunked" ;
		msec:_ChunkSizes = 43200 ;
		msec:_DeflateLevel = 9 ;
		msec:_Shuffle = "true" ;
		msec:_Endianness = "little" ;
	ubyte satID(time) ;
		satID:long_name = "2 digit number identifying the satellite the data is from" ;
		satID:units = "ID" ;
		satID:valid_range = 0., 20. ;
		satID:_Storage = "chunked" ;
		satID:_ChunkSizes = 43200 ;
		satID:_DeflateLevel = 9 ;
		satID:_Shuffle = "true" ;
	ubyte sat_direction(time) ;
		sat_direction:long_name = "satellite direction 0-North/ 1-South" ;
		sat_direction:units = "" ;
		sat_direction:valid_range = 0., 1. ;
		sat_direction:_Storage = "chunked" ;
		sat_direction:_ChunkSizes = 43200 ;
		sat_direction:_DeflateLevel = 9 ;
		sat_direction:_Shuffle = "true" ;
	float alt(time) ;
		alt:long_name = "altitude of the satellite" ;
		alt:units = "km" ;
		alt:valid_range = 800., 1000. ;
		alt:_Storage = "chunked" ;
		alt:_ChunkSizes = 43200 ;
		alt:_DeflateLevel = 9 ;
		alt:_Shuffle = "true" ;
		alt:_FillValue = -1e+31 ;
	float lat(time) ;
		lat:long_name = "latitude of the satellite" ;
		lat:units = "degrees" ;
		lat:valid_range = -90., 90. ;
		lat:_Storage = "chunked" ;
		lat:_ChunkSizes = 43200 ;
		lat:_DeflateLevel = 9 ;
		lat:_Shuffle = "true" ;
		lat:_FillValue = -1e+31 ;
	float lon(time) ;
		lon:long_name = "longitude of the satellite" ;
		lon:units = "degrees" ;
		lon:valid_range = 0., 360. ;
		lon:_Storage = "chunked" ;
		lon:_ChunkSizes = 43200 ;
		lon:_DeflateLevel = 9 ;
		lon:_Shuffle = "true" ;
		lon:_FillValue = -1e+31 ;
	float mep_pro_tel0_flux_p1(time) ;
		mep_pro_tel0_flux_p1:long_name = "MEPED proton flux ~39 keV  0 deg telescope" ;
		mep_pro_tel0_flux_p1:units = "#/cm2-s-str-keV" ;
		mep_pro_tel0_flux_p1:valid_min = 0. ;
		mep_pro_tel0_flux_p1:_Storage = "chunked" ;
		mep_pro_tel0_flux_p1:_ChunkSizes = 43200 ;
		mep_pro_tel0_flux_p1:_DeflateLevel = 9 ;
		mep_pro_tel0_flux_p1:_Shuffle = "true" ;
		mep_pro_tel0_flux_p1:_FillValue = -1e+31 ;
	float mep_pro_tel0_flux_p2(time) ;
		mep_pro_tel0_flux_p2:long_name = "MEPED proton flux ~ 115keV  0 deg telescope" ;
		mep_pro_tel0_flux_p2:units = "#/cm2-s-str-keV" ;
		mep_pro_tel0_flux_p2:valid_min = 0. ;
		mep_pro_tel0_flux_p2:_Storage = "chunked" ;
		mep_pro_tel0_flux_p2:_ChunkSizes = 43200 ;
		mep_pro_tel0_flux_p2:_DeflateLevel = 9 ;
		mep_pro_tel0_flux_p2:_Shuffle = "true" ;
		mep_pro_tel0_flux_p2:_FillValue = -1e+31 ;
	float mep_pro_tel0_flux_p3(time) ;
		mep_pro_tel0_flux_p3:long_name = "MEPED proton flux ~332 keV 0 deg telescope" ;
		mep_pro_tel0_flux_p3:units = "#/cm2-s-str-keV" ;
		mep_pro_tel0_flux_p3:valid_min = 0. ;
		mep_pro_tel0_flux_p3:_Storage = "chunked" ;
		mep_pro_tel0_flux_p3:_ChunkSizes = 43200 ;
		mep_pro_tel0_flux_p3:_DeflateLevel = 9 ;
		mep_pro_tel0_flux_p3:_Shuffle = "true" ;
		mep_pro_tel0_flux_p3:_FillValue = -1e+31 ;
	float mep_pro_tel0_flux_p4(time) ;
		mep_pro_tel0_flux_p4:long_name = "MEPED proton flux ~1105 keV 0 deg telescope" ;
		mep_pro_tel0_flux_p4:units = "#/cm2-s-str-keV" ;
		mep_pro_tel0_flux_p4:valid_min = 0. ;
		mep_pro_tel0_flux_p4:_Storage = "chunked" ;
		mep_pro_tel0_flux_p4:_ChunkSizes = 43200 ;
		mep_pro_tel0_flux_p4:_DeflateLevel = 9 ;
		mep_pro_tel0_flux_p4:_Shuffle = "true" ;
		mep_pro_tel0_flux_p4:_FillValue = -1e+31 ;
	float mep_pro_tel0_flux_p5(time) ;
		mep_pro_tel0_flux_p5:long_name = "MEPED proton flux ~2723 keV 0 deg telescope" ;
		mep_pro_tel0_flux_p5:units = "#/cm2-s-str-keV" ;
		mep_pro_tel0_flux_p5:valid_min = 0. ;
		mep_pro_tel0_flux_p5:_Storage = "chunked" ;
		mep_pro_tel0_flux_p5:_ChunkSizes = 43200 ;
		mep_pro_tel0_flux_p5:_DeflateLevel = 9 ;
		mep_pro_tel0_flux_p5:_Shuffle = "true" ;
		mep_pro_tel0_flux_p5:_FillValue = -1e+31 ;
	float mep_pro_tel0_flux_p6(time) ;
		mep_pro_tel0_flux_p6:long_name = "MEPED proton flux ~6174 keV 0 deg telescope" ;
		mep_pro_tel0_flux_p6:units = "#/cm2-s-str" ;
		mep_pro_tel0_flux_p6:valid_min = 0. ;
		mep_pro_tel0_flux_p6:_Storage = "chunked" ;
		mep_pro_tel0_flux_p6:_ChunkSizes = 43200 ;
		mep_pro_tel0_flux_p6:_DeflateLevel = 9 ;
		mep_pro_tel0_flux_p6:_Shuffle = "true" ;
		mep_pro_tel0_flux_p6:_FillValue = -1e+31 ;
	ushort mep_pro_tel0_flux_p1_err(time) ;
		mep_pro_tel0_flux_p1_err:long_name = "MEPED proton flux percent error ~39 keV  0 deg telescope" ;
		mep_pro_tel0_flux_p1_err:units = "#/cm2-s-str-keV" ;
		mep_pro_tel0_flux_p1_err:valid_min = 0. ;
		mep_pro_tel0_flux_p1_err:_Storage = "chunked" ;
		mep_pro_tel0_flux_p1_err:_ChunkSizes = 43200 ;
		mep_pro_tel0_flux_p1_err:_DeflateLevel = 9 ;
		mep_pro_tel0_flux_p1_err:_Shuffle = "true" ;
		mep_pro_tel0_flux_p1_err:_Endianness = "little" ;
		mep_pro_tel0_flux_p1_err:_FillValue = 65535 ;
	ushort mep_pro_tel0_flux_p2_err(time) ;
		mep_pro_tel0_flux_p2_err:long_name = "MEPED proton flux percent error ~115 keV  0 deg telescope" ;
		mep_pro_tel0_flux_p2_err:units = "#/cm2-s-str-keV" ;
		mep_pro_tel0_flux_p2_err:valid_min = 0. ;
		mep_pro_tel0_flux_p2_err:_Storage = "chunked" ;
		mep_pro_tel0_flux_p2_err:_ChunkSizes = 43200 ;
		mep_pro_tel0_flux_p2_err:_DeflateLevel = 9 ;
		mep_pro_tel0_flux_p2_err:_Shuffle = "true" ;
		mep_pro_tel0_flux_p2_err:_Endianness = "little" ;
		mep_pro_tel0_flux_p2_err:_FillValue = 65535 ;
	ushort mep_pro_tel0_flux_p3_err(time) ;
		mep_pro_tel0_flux_p3_err:long_name = "MEPED proton flux percent error ~332 keV 0 deg telescope" ;
		mep_pro_tel0_flux_p3_err:units = "#/cm2-s-str-keV" ;
		mep_pro_tel0_flux_p3_err:valid_min = 0. ;
		mep_pro_tel0_flux_p3_err:_Storage = "chunked" ;
		mep_pro_tel0_flux_p3_err:_ChunkSizes = 43200 ;
		mep_pro_tel0_flux_p3_err:_DeflateLevel = 9 ;
		mep_pro_tel0_flux_p3_err:_Shuffle = "true" ;
		mep_pro_tel0_flux_p3_err:_Endianness = "little" ;
		mep_pro_tel0_flux_p3_err:_FillValue = 65535 ;
	ushort mep_pro_tel0_flux_p4_err(time) ;
		mep_pro_tel0_flux_p4_err:long_name = "MEPED proton flux percent error ~ 1105keV 0 deg telescope" ;
		mep_pro_tel0_flux_p4_err:units = "#/cm2-s-str-keV" ;
		mep_pro_tel0_flux_p4_err:valid_min = 0. ;
		mep_pro_tel0_flux_p4_err:_Storage = "chunked" ;
		mep_pro_tel0_flux_p4_err:_ChunkSizes = 43200 ;
		mep_pro_tel0_flux_p4_err:_DeflateLevel = 9 ;
		mep_pro_tel0_flux_p4_err:_Shuffle = "true" ;
		mep_pro_tel0_flux_p4_err:_Endianness = "little" ;
		mep_pro_tel0_flux_p4_err:_FillValue = 65535 ;
	ushort mep_pro_tel0_flux_p5_err(time) ;
		mep_pro_tel0_flux_p5_err:long_name = "MEPED proton flux percent error ~2723 keV 0 deg telescope" ;
		mep_pro_tel0_flux_p5_err:units = "#/cm2-s-str-keV" ;
		mep_pro_tel0_flux_p5_err:valid_min = 0. ;
		mep_pro_tel0_flux_p5_err:_Storage = "chunked" ;
		mep_pro_tel0_flux_p5_err:_ChunkSizes = 43200 ;
		mep_pro_tel0_flux_p5_err:_DeflateLevel = 9 ;
		mep_pro_tel0_flux_p5_err:_Shuffle = "true" ;
		mep_pro_tel0_flux_p5_err:_Endianness = "little" ;
		mep_pro_tel0_flux_p5_err:_FillValue = 65535 ;
	ushort mep_pro_tel0_flux_p6_err(time) ;
		mep_pro_tel0_flux_p6_err:long_name = "MEPED proton flux percent error ~6174 keV 0 deg telescope" ;
		mep_pro_tel0_flux_p6_err:units = "#/cm2-s-str" ;
		mep_pro_tel0_flux_p6_err:valid_min = 0. ;
		mep_pro_tel0_flux_p6_err:_Storage = "chunked" ;
		mep_pro_tel0_flux_p6_err:_ChunkSizes = 43200 ;
		mep_pro_tel0_flux_p6_err:_DeflateLevel = 9 ;
		mep_pro_tel0_flux_p6_err:_Shuffle = "true" ;
		mep_pro_tel0_flux_p6_err:_Endianness = "little" ;
		mep_pro_tel0_flux_p6_err:_FillValue = 65535 ;
	float mep_pro_tel90_flux_p1(time) ;
		mep_pro_tel90_flux_p1:long_name = "MEPED proton flux ~39 keV 90 deg telescope" ;
		mep_pro_tel90_flux_p1:units = "#/cm2-s-str-keV" ;
		mep_pro_tel90_flux_p1:valid_min = 0. ;
		mep_pro_tel90_flux_p1:_Storage = "chunked" ;
		mep_pro_tel90_flux_p1:_ChunkSizes = 43200 ;
		mep_pro_tel90_flux_p1:_DeflateLevel = 9 ;
		mep_pro_tel90_flux_p1:_Shuffle = "true" ;
		mep_pro_tel90_flux_p1:_FillValue = -1e+31 ;
	float mep_pro_tel90_flux_p2(time) ;
		mep_pro_tel90_flux_p2:long_name = "MEPED proton flux ~115 keV 90 deg telescope" ;
		mep_pro_tel90_flux_p2:units = "#/cm2-s-str-keV" ;
		mep_pro_tel90_flux_p2:valid_min = 0. ;
		mep_pro_tel90_flux_p2:_Storage = "chunked" ;
		mep_pro_tel90_flux_p2:_ChunkSizes = 43200 ;
		mep_pro_tel90_flux_p2:_DeflateLevel = 9 ;
		mep_pro_tel90_flux_p2:_Shuffle = "true" ;
		mep_pro_tel90_flux_p2:_FillValue = -1e+31 ;
	float mep_pro_tel90_flux_p3(time) ;
		mep_pro_tel90_flux_p3:long_name = "MEPED proton flux ~332 keV 90 deg telescope" ;
		mep_pro_tel90_flux_p3:units = "#/cm2-s-str-keV" ;
		mep_pro_tel90_flux_p3:valid_min = 0. ;
		mep_pro_tel90_flux_p3:_Storage = "chunked" ;
		mep_pro_tel90_flux_p3:_ChunkSizes = 43200 ;
		mep_pro_tel90_flux_p3:_DeflateLevel = 9 ;
		mep_pro_tel90_flux_p3:_Shuffle = "true" ;
		mep_pro_tel90_flux_p3:_FillValue = -1e+31 ;
	float mep_pro_tel90_flux_p4(time) ;
		mep_pro_tel90_flux_p4:long_name = "MEPED proton flux ~1105 keV 90 deg telescope" ;
		mep_pro_tel90_flux_p4:units = "#/cm2-s-str-keV" ;
		mep_pro_tel90_flux_p4:valid_min = 0. ;
		mep_pro_tel90_flux_p4:_Storage = "chunked" ;
		mep_pro_tel90_flux_p4:_ChunkSizes = 43200 ;
		mep_pro_tel90_flux_p4:_DeflateLevel = 9 ;
		mep_pro_tel90_flux_p4:_Shuffle = "true" ;
		mep_pro_tel90_flux_p4:_FillValue = -1e+31 ;
	float mep_pro_tel90_flux_p5(time) ;
		mep_pro_tel90_flux_p5:long_name = "MEPED proton flux ~2723 keV 90 deg telescope" ;
		mep_pro_tel90_flux_p5:units = "#/cm2-s-str-keV" ;
		mep_pro_tel90_flux_p5:valid_min = 0. ;
		mep_pro_tel90_flux_p5:_Storage = "chunked" ;
		mep_pro_tel90_flux_p5:_ChunkSizes = 43200 ;
		mep_pro_tel90_flux_p5:_DeflateLevel = 9 ;
		mep_pro_tel90_flux_p5:_Shuffle = "true" ;
		mep_pro_tel90_flux_p5:_FillValue = -1e+31 ;
	float mep_pro_tel90_flux_p6(time) ;
		mep_pro_tel90_flux_p6:long_name = "MEPED proton flux ~6174 keV 90 deg telescope" ;
		mep_pro_tel90_flux_p6:units = "#/cm2-s-str" ;
		mep_pro_tel90_flux_p6:valid_min = 0. ;
		mep_pro_tel90_flux_p6:_Storage = "chunked" ;
		mep_pro_tel90_flux_p6:_ChunkSizes = 43200 ;
		mep_pro_tel90_flux_p6:_DeflateLevel = 9 ;
		mep_pro_tel90_flux_p6:_Shuffle = "true" ;
		mep_pro_tel90_flux_p6:_FillValue = -1e+31 ;
	short mep_pro_tel90_flux_p1_err(time) ;
		mep_pro_tel90_flux_p1_err:long_name = "MEPED proton flux percent error ~39 keV 90 deg telescope" ;
		mep_pro_tel90_flux_p1_err:units = "#/cm2-s-str-keV" ;
		mep_pro_tel90_flux_p1_err:valid_min = 0. ;
		mep_pro_tel90_flux_p1_err:_Storage = "chunked" ;
		mep_pro_tel90_flux_p1_err:_ChunkSizes = 43200 ;
		mep_pro_tel90_flux_p1_err:_DeflateLevel = 9 ;
		mep_pro_tel90_flux_p1_err:_Shuffle = "true" ;
		mep_pro_tel90_flux_p1_err:_Endianness = "little" ;
		mep_pro_tel90_flux_p1_err:_FillValue = -32767 ;
	short mep_pro_tel90_flux_p2_err(time) ;
		mep_pro_tel90_flux_p2_err:long_name = "MEPED proton flux percent error ~115 keV 90 deg telescope" ;
		mep_pro_tel90_flux_p2_err:units = "#/cm2-s-str-keV" ;
		mep_pro_tel90_flux_p2_err:valid_min = 0. ;
		mep_pro_tel90_flux_p2_err:_Storage = "chunked" ;
		mep_pro_tel90_flux_p2_err:_ChunkSizes = 43200 ;
		mep_pro_tel90_flux_p2_err:_DeflateLevel = 9 ;
		mep_pro_tel90_flux_p2_err:_Shuffle = "true" ;
		mep_pro_tel90_flux_p2_err:_Endianness = "little" ;
		mep_pro_tel90_flux_p2_err:_FillValue = -32767 ;
	short mep_pro_tel90_flux_p3_err(time) ;
		mep_pro_tel90_flux_p3_err:long_name = "MEPED proton flux percent error ~332 keV 90 deg telescope" ;
		mep_pro_tel90_flux_p3_err:units = "#/cm2-s-str-keV" ;
		mep_pro_tel90_flux_p3_err:valid_min = 0. ;
		mep_pro_tel90_flux_p3_err:_Storage = "chunked" ;
		mep_pro_tel90_flux_p3_err:_ChunkSizes = 43200 ;
		mep_pro_tel90_flux_p3_err:_DeflateLevel = 9 ;
		mep_pro_tel90_flux_p3_err:_Shuffle = "true" ;
		mep_pro_tel90_flux_p3_err:_Endianness = "little" ;
		mep_pro_tel90_flux_p3_err:_FillValue = -32767 ;
	short mep_pro_tel90_flux_p4_err(time) ;
		mep_pro_tel90_flux_p4_err:long_name = "MEPED proton flux percent error ~1105 keV 90 deg telescope" ;
		mep_pro_tel90_flux_p4_err:units = "#/cm2-s-str-keV" ;
		mep_pro_tel90_flux_p4_err:valid_min = 0. ;
		mep_pro_tel90_flux_p4_err:_Storage = "chunked" ;
		mep_pro_tel90_flux_p4_err:_ChunkSizes = 43200 ;
		mep_pro_tel90_flux_p4_err:_DeflateLevel = 9 ;
		mep_pro_tel90_flux_p4_err:_Shuffle = "true" ;
		mep_pro_tel90_flux_p4_err:_Endianness = "little" ;
		mep_pro_tel90_flux_p4_err:_FillValue = -32767 ;
	short mep_pro_tel90_flux_p5_err(time) ;
		mep_pro_tel90_flux_p5_err:long_name = "MEPED proton flux percent error ~2723 keV 90 deg telescope" ;
		mep_pro_tel90_flux_p5_err:units = "#/cm2-s-str-keV" ;
		mep_pro_tel90_flux_p5_err:valid_min = 0. ;
		mep_pro_tel90_flux_p5_err:_Storage = "chunked" ;
		mep_pro_tel90_flux_p5_err:_ChunkSizes = 43200 ;
		mep_pro_tel90_flux_p5_err:_DeflateLevel = 9 ;
		mep_pro_tel90_flux_p5_err:_Shuffle = "true" ;
		mep_pro_tel90_flux_p5_err:_Endianness = "little" ;
		mep_pro_tel90_flux_p5_err:_FillValue = -32767 ;
	short mep_pro_tel90_flux_p6_err(time) ;
		mep_pro_tel90_flux_p6_err:long_name = "MEPED proton flux percent error ~6174 keV 90 deg telescope" ;
		mep_pro_tel90_flux_p6_err:units = "#/cm2-s-str" ;
		mep_pro_tel90_flux_p6_err:valid_min = 0. ;
		mep_pro_tel90_flux_p6_err:_Storage = "chunked" ;
		mep_pro_tel90_flux_p6_err:_ChunkSizes = 43200 ;
		mep_pro_tel90_flux_p6_err:_DeflateLevel = 9 ;
		mep_pro_tel90_flux_p6_err:_Shuffle = "true" ;
		mep_pro_tel90_flux_p6_err:_Endianness = "little" ;
		mep_pro_tel90_flux_p6_err:_FillValue = -32767 ;
	float mep_ele_tel0_flux_e1(time) ;
		mep_ele_tel0_flux_e1:long_name = "MEPED electron flux >40 keV 0 deg telescope" ;
		mep_ele_tel0_flux_e1:units = "#/cm2-s-str" ;
		mep_ele_tel0_flux_e1:valid_min = 0. ;
		mep_ele_tel0_flux_e1:_Storage = "chunked" ;
		mep_ele_tel0_flux_e1:_ChunkSizes = 43200 ;
		mep_ele_tel0_flux_e1:_DeflateLevel = 9 ;
		mep_ele_tel0_flux_e1:_Shuffle = "true" ;
		mep_ele_tel0_flux_e1:_FillValue = -1e+31 ;
	float mep_ele_tel0_flux_e2(time) ;
		mep_ele_tel0_flux_e2:long_name = "MEPED electron flux >130 keV 0 deg telescope" ;
		mep_ele_tel0_flux_e2:units = "#/cm2-s-str" ;
		mep_ele_tel0_flux_e2:valid_min = 0. ;
		mep_ele_tel0_flux_e2:_Storage = "chunked" ;
		mep_ele_tel0_flux_e2:_ChunkSizes = 43200 ;
		mep_ele_tel0_flux_e2:_DeflateLevel = 9 ;
		mep_ele_tel0_flux_e2:_Shuffle = "true" ;
		mep_ele_tel0_flux_e2:_FillValue = -1e+31 ;
	float mep_ele_tel0_flux_e3(time) ;
		mep_ele_tel0_flux_e3:long_name = "MEPED electron flux >287 keV 0 deg telescope" ;
		mep_ele_tel0_flux_e3:units = "#/cm2-s-str" ;
		mep_ele_tel0_flux_e3:valid_min = 0. ;
		mep_ele_tel0_flux_e3:_Storage = "chunked" ;
		mep_ele_tel0_flux_e3:_ChunkSizes = 43200 ;
		mep_ele_tel0_flux_e3:_DeflateLevel = 9 ;
		mep_ele_tel0_flux_e3:_Shuffle = "true" ;
		mep_ele_tel0_flux_e3:_FillValue = -1e+31 ;
	float mep_ele_tel0_flux_e4(time) ;
		mep_ele_tel0_flux_e4:long_name = "MEPED electron flux >612 keV 0 deg telescope" ;
		mep_ele_tel0_flux_e4:units = "#/cm2-s-str" ;
		mep_ele_tel0_flux_e4:valid_min = 0. ;
		mep_ele_tel0_flux_e4:_Storage = "chunked" ;
		mep_ele_tel0_flux_e4:_ChunkSizes = 43200 ;
		mep_ele_tel0_flux_e4:_DeflateLevel = 9 ;
		mep_ele_tel0_flux_e4:_Shuffle = "true" ;
		mep_ele_tel0_flux_e4:_FillValue = -1e+31 ;
	short mep_ele_tel0_flux_e1_err(time) ;
		mep_ele_tel0_flux_e1_err:long_name = "MEPED electron flux percent error >40 keV 0 deg telescope" ;
		mep_ele_tel0_flux_e1_err:units = "#/cm2-s-str" ;
		mep_ele_tel0_flux_e1_err:valid_min = 0. ;
		mep_ele_tel0_flux_e1_err:_Storage = "chunked" ;
		mep_ele_tel0_flux_e1_err:_ChunkSizes = 43200 ;
		mep_ele_tel0_flux_e1_err:_DeflateLevel = 9 ;
		mep_ele_tel0_flux_e1_err:_Shuffle = "true" ;
		mep_ele_tel0_flux_e1_err:_Endianness = "little" ;
		mep_ele_tel0_flux_e1_err:_FillValue = -32767 ;
	short mep_ele_tel0_flux_e2_err(time) ;
		mep_ele_tel0_flux_e2_err:long_name = "MEPED electron flux percent error >130 keV 0 deg telescope" ;
		mep_ele_tel0_flux_e2_err:units = "#/cm2-s-str" ;
		mep_ele_tel0_flux_e2_err:valid_min = 0. ;
		mep_ele_tel0_flux_e2_err:_Storage = "chunked" ;
		mep_ele_tel0_flux_e2_err:_ChunkSizes = 43200 ;
		mep_ele_tel0_flux_e2_err:_DeflateLevel = 9 ;
		mep_ele_tel0_flux_e2_err:_Shuffle = "true" ;
		mep_ele_tel0_flux_e2_err:_Endianness = "little" ;
		mep_ele_tel0_flux_e2_err:_FillValue = -32767 ;
	short mep_ele_tel0_flux_e3_err(time) ;
		mep_ele_tel0_flux_e3_err:long_name = "MEPED electron flux percent error >287 keV 0 deg telescope" ;
		mep_ele_tel0_flux_e3_err:units = "#/cm2-s-str" ;
		mep_ele_tel0_flux_e3_err:valid_min = 0. ;
		mep_ele_tel0_flux_e3_err:_Storage = "chunked" ;
		mep_ele_tel0_flux_e3_err:_ChunkSizes = 43200 ;
		mep_ele_tel0_flux_e3_err:_DeflateLevel = 9 ;
		mep_ele_tel0_flux_e3_err:_Shuffle = "true" ;
		mep_ele_tel0_flux_e3_err:_Endianness = "little" ;
		mep_ele_tel0_flux_e3_err:_FillValue = -32767 ;
	short mep_ele_tel0_flux_e4_err(time) ;
		mep_ele_tel0_flux_e4_err:long_name = "MEPED electron flux percent error >612 keV 0 deg telescope" ;
		mep_ele_tel0_flux_e4_err:units = "#/cm2-s-str" ;
		mep_ele_tel0_flux_e4_err:valid_min = 0. ;
		mep_ele_tel0_flux_e4_err:_Storage = "chunked" ;
		mep_ele_tel0_flux_e4_err:_ChunkSizes = 43200 ;
		mep_ele_tel0_flux_e4_err:_DeflateLevel = 9 ;
		mep_ele_tel0_flux_e4_err:_Shuffle = "true" ;
		mep_ele_tel0_flux_e4_err:_Endianness = "little" ;
		mep_ele_tel0_flux_e4_err:_FillValue = -32767 ;
	float mep_ele_tel90_flux_e1(time) ;
		mep_ele_tel90_flux_e1:long_name = "MEPED electron flux >40 keV 90 deg telescope" ;
		mep_ele_tel90_flux_e1:units = "#/cm2-s-str" ;
		mep_ele_tel90_flux_e1:valid_min = 0. ;
		mep_ele_tel90_flux_e1:_Storage = "chunked" ;
		mep_ele_tel90_flux_e1:_ChunkSizes = 43200 ;
		mep_ele_tel90_flux_e1:_DeflateLevel = 9 ;
		mep_ele_tel90_flux_e1:_Shuffle = "true" ;
		mep_ele_tel90_flux_e1:_FillValue = -1e+31 ;
	float mep_ele_tel90_flux_e2(time) ;
		mep_ele_tel90_flux_e2:long_name = "MEPED electron flux >130 keV 90 deg telescope" ;
		mep_ele_tel90_flux_e2:units = "#/cm2-s-str" ;
		mep_ele_tel90_flux_e2:valid_min = 0. ;
		mep_ele_tel90_flux_e2:_Storage = "chunked" ;
		mep_ele_tel90_flux_e2:_ChunkSizes = 43200 ;
		mep_ele_tel90_flux_e2:_DeflateLevel = 9 ;
		mep_ele_tel90_flux_e2:_Shuffle = "true" ;
		mep_ele_tel90_flux_e2:_FillValue = -1e+31 ;
	float mep_ele_tel90_flux_e3(time) ;
		mep_ele_tel90_flux_e3:long_name = "MEPED electron flux >287 keV 90 deg telescope" ;
		mep_ele_tel90_flux_e3:units = "#/cm2-s-str" ;
		mep_ele_tel90_flux_e3:valid_min = 0. ;
		mep_ele_tel90_flux_e3:_Storage = "chunked" ;
		mep_ele_tel90_flux_e3:_ChunkSizes = 43200 ;
		mep_ele_tel90_flux_e3:_DeflateLevel = 9 ;
		mep_ele_tel90_flux_e3:_Shuffle = "true" ;
		mep_ele_tel90_flux_e3:_FillValue = -1e+31 ;
	float mep_ele_tel90_flux_e4(time) ;
		mep_ele_tel90_flux_e4:long_name = "MEPED electron flux >6174 keV 90 deg telescope" ;
		mep_ele_tel90_flux_e4:units = "#/cm2-s-str" ;
		mep_ele_tel90_flux_e4:valid_min = 0. ;
		mep_ele_tel90_flux_e4:_Storage = "chunked" ;
		mep_ele_tel90_flux_e4:_ChunkSizes = 43200 ;
		mep_ele_tel90_flux_e4:_DeflateLevel = 9 ;
		mep_ele_tel90_flux_e4:_Shuffle = "true" ;
		mep_ele_tel90_flux_e4:_FillValue = -1e+31 ;
	short mep_ele_tel90_flux_e1_err(time) ;
		mep_ele_tel90_flux_e1_err:long_name = "MEPED electron flux percent error >40 keV 90 deg telescope" ;
		mep_ele_tel90_flux_e1_err:units = "#/cm2-s-str" ;
		mep_ele_tel90_flux_e1_err:valid_min = 0. ;
		mep_ele_tel90_flux_e1_err:_Storage = "chunked" ;
		mep_ele_tel90_flux_e1_err:_ChunkSizes = 43200 ;
		mep_ele_tel90_flux_e1_err:_DeflateLevel = 9 ;
		mep_ele_tel90_flux_e1_err:_Shuffle = "true" ;
		mep_ele_tel90_flux_e1_err:_Endianness = "little" ;
		mep_ele_tel90_flux_e1_err:_FillValue = -32767 ;
	short mep_ele_tel90_flux_e2_err(time) ;
		mep_ele_tel90_flux_e2_err:long_name = "MEPED electron flux percent error >130 keV 90 deg telescope" ;
		mep_ele_tel90_flux_e2_err:units = "#/cm2-s-str" ;
		mep_ele_tel90_flux_e2_err:valid_min = 0. ;
		mep_ele_tel90_flux_e2_err:_Storage = "chunked" ;
		mep_ele_tel90_flux_e2_err:_ChunkSizes = 43200 ;
		mep_ele_tel90_flux_e2_err:_DeflateLevel = 9 ;
		mep_ele_tel90_flux_e2_err:_Shuffle = "true" ;
		mep_ele_tel90_flux_e2_err:_Endianness = "little" ;
		mep_ele_tel90_flux_e2_err:_FillValue = -32767 ;
	short mep_ele_tel90_flux_e3_err(time) ;
		mep_ele_tel90_flux_e3_err:long_name = "MEPED electron flux percent error >287 keV 90 deg telescope" ;
		mep_ele_tel90_flux_e3_err:units = "#/cm2-s-str" ;
		mep_ele_tel90_flux_e3_err:valid_min = 0. ;
		mep_ele_tel90_flux_e3_err:_Storage = "chunked" ;
		mep_ele_tel90_flux_e3_err:_ChunkSizes = 43200 ;
		mep_ele_tel90_flux_e3_err:_DeflateLevel = 9 ;
		mep_ele_tel90_flux_e3_err:_Shuffle = "true" ;
		mep_ele_tel90_flux_e3_err:_Endianness = "little" ;
		mep_ele_tel90_flux_e3_err:_FillValue = -32767 ;
	short mep_ele_tel90_flux_e4_err(time) ;
		mep_ele_tel90_flux_e4_err:long_name = "MEPED electron flux percent error >6174 keV 90 deg telescope" ;
		mep_ele_tel90_flux_e4_err:units = "#/cm2-s-str" ;
		mep_ele_tel90_flux_e4_err:valid_min = 0. ;
		mep_ele_tel90_flux_e4_err:_Storage = "chunked" ;
		mep_ele_tel90_flux_e4_err:_ChunkSizes = 43200 ;
		mep_ele_tel90_flux_e4_err:_DeflateLevel = 9 ;
		mep_ele_tel90_flux_e4_err:_Shuffle = "true" ;
		mep_ele_tel90_flux_e4_err:_Endianness = "little" ;
		mep_ele_tel90_flux_e4_err:_FillValue = -32767 ;
	float mep_omni_flux_p1(time) ;
		mep_omni_flux_p1:long_name = "MEPED proton differential flux at 25 MeV omnidirection telescope" ;
		mep_omni_flux_p1:units = "#/cm2-s-str-MeV" ;
		mep_omni_flux_p1:valid_min = 0. ;
		mep_omni_flux_p1:_Storage = "chunked" ;
		mep_omni_flux_p1:_ChunkSizes = 43200 ;
		mep_omni_flux_p1:_DeflateLevel = 9 ;
		mep_omni_flux_p1:_Shuffle = "true" ;
		mep_omni_flux_p1:_FillValue = -1e+31 ;
	float mep_omni_flux_p2(time) ;
		mep_omni_flux_p2:long_name = "MEPED proton differential flux at 50 MeV omnidirection telescope" ;
		mep_omni_flux_p2:units = "#/cm2-s-str-MeV" ;
		mep_omni_flux_p2:valid_min = 0. ;
		mep_omni_flux_p2:_Storage = "chunked" ;
		mep_omni_flux_p2:_ChunkSizes = 43200 ;
		mep_omni_flux_p2:_DeflateLevel = 9 ;
		mep_omni_flux_p2:_Shuffle = "true" ;
		mep_omni_flux_p2:_FillValue = -1e+31 ;
	float mep_omni_flux_p3(time) ;
		mep_omni_flux_p3:long_name = "MEPED proton differential flux at 100 MeV omnidirection telescope" ;
		mep_omni_flux_p3:units = "#/cm2-s-str-MeV" ;
		mep_omni_flux_p3:valid_min = 0. ;
		mep_omni_flux_p3:_Storage = "chunked" ;
		mep_omni_flux_p3:_ChunkSizes = 43200 ;
		mep_omni_flux_p3:_DeflateLevel = 9 ;
		mep_omni_flux_p3:_Shuffle = "true" ;
		mep_omni_flux_p3:_FillValue = -1e+31 ;
	byte mep_omni_flux_flag_fit(time) ;
		mep_omni_flux_flag_fit:long_name = "MEPED omni fit flag" ;
		mep_omni_flux_flag_fit:units = "flag" ;
		mep_omni_flux_flag_fit:valid_range = -1., 2. ;
		mep_omni_flux_flag_fit:_Storage = "chunked" ;
		mep_omni_flux_flag_fit:_ChunkSizes = 43200 ;
		mep_omni_flux_flag_fit:_DeflateLevel = 9 ;
		mep_omni_flux_flag_fit:_Shuffle = "true" ;
	byte mep_omni_flux_flag_iter_lim(time) ;
		mep_omni_flux_flag_iter_lim:long_name = "MEPED omni flag for fit iteration limit" ;
		mep_omni_flux_flag_iter_lim:units = "true/false" ;
		mep_omni_flux_flag_iter_lim:valid_range = 0., 1. ;
		mep_omni_flux_flag_iter_lim:_Storage = "chunked" ;
		mep_omni_flux_flag_iter_lim:_ChunkSizes = 43200 ;
		mep_omni_flux_flag_iter_lim:_DeflateLevel = 9 ;
		mep_omni_flux_flag_iter_lim:_Shuffle = "true" ;
	float mep_omni_gamma_p1(time) ;
		mep_omni_gamma_p1:long_name = "gamma derived for p1 energy band" ;
		mep_omni_gamma_p1:units = "" ;
		mep_omni_gamma_p1:_Storage = "chunked" ;
		mep_omni_gamma_p1:_ChunkSizes = 43200 ;
		mep_omni_gamma_p1:_DeflateLevel = 9 ;
		mep_omni_gamma_p1:_Shuffle = "true" ;
		mep_omni_gamma_p1:_FillValue = -1e+31 ;
	float mep_omni_gamma_p2(time) ;
		mep_omni_gamma_p2:long_name = "gamma derived for p2 energy band" ;
		mep_omni_gamma_p2:units = "" ;
		mep_omni_gamma_p2:_Storage = "chunked" ;
		mep_omni_gamma_p2:_ChunkSizes = 43200 ;
		mep_omni_gamma_p2:_DeflateLevel = 9 ;
		mep_omni_gamma_p2:_Shuffle = "true" ;
		mep_omni_gamma_p2:_FillValue = -1e+31 ;
	float mep_omni_gamma_p3(time) ;
		mep_omni_gamma_p3:long_name = "gamma derived for p3 energy band" ;
		mep_omni_gamma_p3:units = "" ;
		mep_omni_gamma_p3:_Storage = "chunked" ;
		mep_omni_gamma_p3:_ChunkSizes = 43200 ;
		mep_omni_gamma_p3:_DeflateLevel = 9 ;
		mep_omni_gamma_p3:_Shuffle = "true" ;
		mep_omni_gamma_p3:_FillValue = -1e+31 ;
	float ted_ele_tel0_flux_4(time) ;
		ted_ele_tel0_flux_4:long_name = "TED electron 189 eV 0 deg telescope" ;
		ted_ele_tel0_flux_4:units = "[#/cm2-s-str-eV]" ;
		ted_ele_tel0_flux_4:valid_range = 0., 4000000000. ;
		ted_ele_tel0_flux_4:_Storage = "chunked" ;
		ted_ele_tel0_flux_4:_ChunkSizes = 43200 ;
		ted_ele_tel0_flux_4:_DeflateLevel = 9 ;
		ted_ele_tel0_flux_4:_Shuffle = "true" ;
		ted_ele_tel0_flux_4:_FillValue = -1e+31 ;
	float ted_ele_tel0_flux_8(time) ;
		ted_ele_tel0_flux_8:long_name = "TED electron 844 eV 0 deg telescope" ;
		ted_ele_tel0_flux_8:units = "[#/cm2-s-str-eV]" ;
		ted_ele_tel0_flux_8:valid_range = 0., 4000000000. ;
		ted_ele_tel0_flux_8:_Storage = "chunked" ;
		ted_ele_tel0_flux_8:_ChunkSizes = 43200 ;
		ted_ele_tel0_flux_8:_DeflateLevel = 9 ;
		ted_ele_tel0_flux_8:_Shuffle = "true" ;
		ted_ele_tel0_flux_8:_FillValue = -1e+31 ;
	float ted_ele_tel0_flux_11(time) ;
		ted_ele_tel0_flux_11:long_name = "TED electron 2595 eV 0 deg telescope" ;
		ted_ele_tel0_flux_11:units = "[#/cm2-s-str-eV]" ;
		ted_ele_tel0_flux_11:valid_range = 0., 4000000000. ;
		ted_ele_tel0_flux_11:_Storage = "chunked" ;
		ted_ele_tel0_flux_11:_ChunkSizes = 43200 ;
		ted_ele_tel0_flux_11:_DeflateLevel = 9 ;
		ted_ele_tel0_flux_11:_Shuffle = "true" ;
		ted_ele_tel0_flux_11:_FillValue = -1e+31 ;
	float ted_ele_tel0_flux_14(time) ;
		ted_ele_tel0_flux_14:long_name = "TED electron 7980 eV 0 deg telescope" ;
		ted_ele_tel0_flux_14:units = "[#/cm2-s-str-eV]" ;
		ted_ele_tel0_flux_14:valid_range = 0., 4000000000. ;
		ted_ele_tel0_flux_14:_Storage = "chunked" ;
		ted_ele_tel0_flux_14:_ChunkSizes = 43200 ;
		ted_ele_tel0_flux_14:_DeflateLevel = 9 ;
		ted_ele_tel0_flux_14:_Shuffle = "true" ;
		ted_ele_tel0_flux_14:_FillValue = -1e+31 ;
	float ted_ele_tel30_flux_4(time) ;
		ted_ele_tel30_flux_4:long_name = "TED electron 189 eV 30 deg telescope" ;
		ted_ele_tel30_flux_4:units = "[#/cm2-s-str-eV]" ;
		ted_ele_tel30_flux_4:valid_range = 0., 4000000000. ;
		ted_ele_tel30_flux_4:_Storage = "chunked" ;
		ted_ele_tel30_flux_4:_ChunkSizes = 43200 ;
		ted_ele_tel30_flux_4:_DeflateLevel = 9 ;
		ted_ele_tel30_flux_4:_Shuffle = "true" ;
		ted_ele_tel30_flux_4:_FillValue = -1e+31 ;
	float ted_ele_tel30_flux_8(time) ;
		ted_ele_tel30_flux_8:long_name = "TED electron 844 eV  30 deg telescope" ;
		ted_ele_tel30_flux_8:units = "[#/cm2-s-str-eV]" ;
		ted_ele_tel30_flux_8:valid_range = 0., 4000000000. ;
		ted_ele_tel30_flux_8:_Storage = "chunked" ;
		ted_ele_tel30_flux_8:_ChunkSizes = 43200 ;
		ted_ele_tel30_flux_8:_DeflateLevel = 9 ;
		ted_ele_tel30_flux_8:_Shuffle = "true" ;
		ted_ele_tel30_flux_8:_FillValue = -1e+31 ;
	float ted_ele_tel30_flux_11(time) ;
		ted_ele_tel30_flux_11:long_name = "TED electron 2595 eV 30 deg telescope" ;
		ted_ele_tel30_flux_11:units = "[#/cm2-s-str-eV]" ;
		ted_ele_tel30_flux_11:valid_range = 0., 4000000000. ;
		ted_ele_tel30_flux_11:_Storage = "chunked" ;
		ted_ele_tel30_flux_11:_ChunkSizes = 43200 ;
		ted_ele_tel30_flux_11:_DeflateLevel = 9 ;
		ted_ele_tel30_flux_11:_Shuffle = "true" ;
		ted_ele_tel30_flux_11:_FillValue = -1e+31 ;
	float ted_ele_tel30_flux_14(time) ;
		ted_ele_tel30_flux_14:long_name = "TED electron 7980 30 deg telescope" ;
		ted_ele_tel30_flux_14:units = "[#/cm2-s-str-eV]" ;
		ted_ele_tel30_flux_14:valid_range = 0., 4000000000. ;
		ted_ele_tel30_flux_14:_Storage = "chunked" ;
		ted_ele_tel30_flux_14:_ChunkSizes = 43200 ;
		ted_ele_tel30_flux_14:_DeflateLevel = 9 ;
		ted_ele_tel30_flux_14:_Shuffle = "true" ;
		ted_ele_tel30_flux_14:_FillValue = -1e+31 ;
	float ted_pro_tel0_flux_4(time) ;
		ted_pro_tel0_flux_4:long_name = "TED proton 189 eV 0 deg telescope" ;
		ted_pro_tel0_flux_4:units = "[#/cm2-s-str-eV]" ;
		ted_pro_tel0_flux_4:valid_range = 0., 4000000000. ;
		ted_pro_tel0_flux_4:_Storage = "chunked" ;
		ted_pro_tel0_flux_4:_ChunkSizes = 43200 ;
		ted_pro_tel0_flux_4:_DeflateLevel = 9 ;
		ted_pro_tel0_flux_4:_Shuffle = "true" ;
		ted_pro_tel0_flux_4:_FillValue = -1e+31 ;
	float ted_pro_tel0_flux_8(time) ;
		ted_pro_tel0_flux_8:long_name = "TED proton 844 eV  0 deg telescope" ;
		ted_pro_tel0_flux_8:units = "[#/cm2-s-str-eV]" ;
		ted_pro_tel0_flux_8:valid_range = 0., 4000000000. ;
		ted_pro_tel0_flux_8:_Storage = "chunked" ;
		ted_pro_tel0_flux_8:_ChunkSizes = 43200 ;
		ted_pro_tel0_flux_8:_DeflateLevel = 9 ;
		ted_pro_tel0_flux_8:_Shuffle = "true" ;
		ted_pro_tel0_flux_8:_FillValue = -1e+31 ;
	float ted_pro_tel0_flux_11(time) ;
		ted_pro_tel0_flux_11:long_name = "TED proton 2595 eV 0 deg telescope" ;
		ted_pro_tel0_flux_11:units = "[#/cm2-s-str-eV]" ;
		ted_pro_tel0_flux_11:valid_range = 0., 4000000000. ;
		ted_pro_tel0_flux_11:_Storage = "chunked" ;
		ted_pro_tel0_flux_11:_ChunkSizes = 43200 ;
		ted_pro_tel0_flux_11:_DeflateLevel = 9 ;
		ted_pro_tel0_flux_11:_Shuffle = "true" ;
		ted_pro_tel0_flux_11:_FillValue = -1e+31 ;
	float ted_pro_tel0_flux_14(time) ;
		ted_pro_tel0_flux_14:long_name = "TED proton 7980 0 deg telescope" ;
		ted_pro_tel0_flux_14:units = "[#/cm2-s-str-eV]" ;
		ted_pro_tel0_flux_14:valid_range = 0., 4000000000. ;
		ted_pro_tel0_flux_14:_Storage = "chunked" ;
		ted_pro_tel0_flux_14:_ChunkSizes = 43200 ;
		ted_pro_tel0_flux_14:_DeflateLevel = 9 ;
		ted_pro_tel0_flux_14:_Shuffle = "true" ;
		ted_pro_tel0_flux_14:_FillValue = -1e+31 ;
	float ted_pro_tel30_flux_4(time) ;
		ted_pro_tel30_flux_4:long_name = "TED proton 189 eV 30 deg telescope" ;
		ted_pro_tel30_flux_4:units = "[#/cm2-s-str-eV]" ;
		ted_pro_tel30_flux_4:valid_range = 0., 4000000000. ;
		ted_pro_tel30_flux_4:_Storage = "chunked" ;
		ted_pro_tel30_flux_4:_ChunkSizes = 43200 ;
		ted_pro_tel30_flux_4:_DeflateLevel = 9 ;
		ted_pro_tel30_flux_4:_Shuffle = "true" ;
		ted_pro_tel30_flux_4:_FillValue = -1e+31 ;
	float ted_pro_tel30_flux_8(time) ;
		ted_pro_tel30_flux_8:long_name = "TED proton 844 eV 30 deg telescope" ;
		ted_pro_tel30_flux_8:units = "[#/cm2-s-str-eV]" ;
		ted_pro_tel30_flux_8:valid_range = 0., 4000000000. ;
		ted_pro_tel30_flux_8:_Storage = "chunked" ;
		ted_pro_tel30_flux_8:_ChunkSizes = 43200 ;
		ted_pro_tel30_flux_8:_DeflateLevel = 9 ;
		ted_pro_tel30_flux_8:_Shuffle = "true" ;
		ted_pro_tel30_flux_8:_FillValue = -1e+31 ;
	float ted_pro_tel30_flux_11(time) ;
		ted_pro_tel30_flux_11:long_name = "TED proton 2595 eV 30 deg telescope" ;
		ted_pro_tel30_flux_11:units = "[#/cm2-s-str-eV]" ;
		ted_pro_tel30_flux_11:valid_range = 0., 4000000000. ;
		ted_pro_tel30_flux_11:_Storage = "chunked" ;
		ted_pro_tel30_flux_11:_ChunkSizes = 43200 ;
		ted_pro_tel30_flux_11:_DeflateLevel = 9 ;
		ted_pro_tel30_flux_11:_Shuffle = "true" ;
		ted_pro_tel30_flux_11:_FillValue = -1e+31 ;
	float ted_pro_tel30_flux_14(time) ;
		ted_pro_tel30_flux_14:long_name = "TED proton 7980 eV 30 deg telescope" ;
		ted_pro_tel30_flux_14:units = "[#/cm2-s-str-eV]" ;
		ted_pro_tel30_flux_14:valid_range = 0., 4000000000. ;
		ted_pro_tel30_flux_14:_Storage = "chunked" ;
		ted_pro_tel30_flux_14:_ChunkSizes = 43200 ;
		ted_pro_tel30_flux_14:_DeflateLevel = 9 ;
		ted_pro_tel30_flux_14:_Shuffle = "true" ;
		ted_pro_tel30_flux_14:_FillValue = -1e+31 ;
	float ted_ele_tel0_low_eflux(time) ;
		ted_ele_tel0_low_eflux:long_name = "TED electron (50eV-1 keV) 0 deg telescope energy flux" ;
		ted_ele_tel0_low_eflux:units = "mW/m2-str" ;
		ted_ele_tel0_low_eflux:valid_range = -200., 200. ;
		ted_ele_tel0_low_eflux:_Storage = "chunked" ;
		ted_ele_tel0_low_eflux:_ChunkSizes = 43200 ;
		ted_ele_tel0_low_eflux:_DeflateLevel = 9 ;
		ted_ele_tel0_low_eflux:_Shuffle = "true" ;
		ted_ele_tel0_low_eflux:_FillValue = -1e+31 ;
	float ted_ele_tel30_low_eflux(time) ;
		ted_ele_tel30_low_eflux:long_name = "TED electron (50eV-1 keV) 30 deg telescope energy flux" ;
		ted_ele_tel30_low_eflux:units = "mW/m2-str" ;
		ted_ele_tel30_low_eflux:valid_range = -200., 200. ;
		ted_ele_tel30_low_eflux:_Storage = "chunked" ;
		ted_ele_tel30_low_eflux:_ChunkSizes = 43200 ;
		ted_ele_tel30_low_eflux:_DeflateLevel = 9 ;
		ted_ele_tel30_low_eflux:_Shuffle = "true" ;
		ted_ele_tel30_low_eflux:_FillValue = -1e+31 ;
	float ted_ele_tel0_hi_eflux(time) ;
		ted_ele_tel0_hi_eflux:long_name = "TED electron (1-20 keV) 0 deg telescope energy flux" ;
		ted_ele_tel0_hi_eflux:units = "mW/m2-str" ;
		ted_ele_tel0_hi_eflux:valid_range = -200., 200. ;
		ted_ele_tel0_hi_eflux:_Storage = "chunked" ;
		ted_ele_tel0_hi_eflux:_ChunkSizes = 43200 ;
		ted_ele_tel0_hi_eflux:_DeflateLevel = 9 ;
		ted_ele_tel0_hi_eflux:_Shuffle = "true" ;
		ted_ele_tel0_hi_eflux:_FillValue = -1e+31 ;
	float ted_ele_tel30_hi_eflux(time) ;
		ted_ele_tel30_hi_eflux:long_name = "TED electron (1-20 keV)  30 deg telescope energy flux" ;
		ted_ele_tel30_hi_eflux:units = "mW/m2-str" ;
		ted_ele_tel30_hi_eflux:valid_range = -200., 200. ;
		ted_ele_tel30_hi_eflux:_Storage = "chunked" ;
		ted_ele_tel30_hi_eflux:_ChunkSizes = 43200 ;
		ted_ele_tel30_hi_eflux:_DeflateLevel = 9 ;
		ted_ele_tel30_hi_eflux:_Shuffle = "true" ;
		ted_ele_tel30_hi_eflux:_FillValue = -1e+31 ;
	float ted_pro_tel0_low_eflux(time) ;
		ted_pro_tel0_low_eflux:long_name = "TED proton (50eV-1 keV) 0 deg telescope energy flux" ;
		ted_pro_tel0_low_eflux:units = "mW/m2-str" ;
		ted_pro_tel0_low_eflux:valid_range = -200., 200. ;
		ted_pro_tel0_low_eflux:_Storage = "chunked" ;
		ted_pro_tel0_low_eflux:_ChunkSizes = 43200 ;
		ted_pro_tel0_low_eflux:_DeflateLevel = 9 ;
		ted_pro_tel0_low_eflux:_Shuffle = "true" ;
		ted_pro_tel0_low_eflux:_FillValue = -1e+31 ;
	float ted_pro_tel30_low_eflux(time) ;
		ted_pro_tel30_low_eflux:long_name = "TEDproton (50eV-1 keV) 30 deg telescope energy flux" ;
		ted_pro_tel30_low_eflux:units = "mW/m2-str" ;
		ted_pro_tel30_low_eflux:valid_range = -200., 200. ;
		ted_pro_tel30_low_eflux:_Storage = "chunked" ;
		ted_pro_tel30_low_eflux:_ChunkSizes = 43200 ;
		ted_pro_tel30_low_eflux:_DeflateLevel = 9 ;
		ted_pro_tel30_low_eflux:_Shuffle = "true" ;
		ted_pro_tel30_low_eflux:_FillValue = -1e+31 ;
	float ted_pro_tel0_hi_eflux(time) ;
		ted_pro_tel0_hi_eflux:long_name = "TED proton (1-20 keV)  0 deg telescope energy flux" ;
		ted_pro_tel0_hi_eflux:units = "mW/m2-str" ;
		ted_pro_tel0_hi_eflux:valid_range = -200., 200. ;
		ted_pro_tel0_hi_eflux:_Storage = "chunked" ;
		ted_pro_tel0_hi_eflux:_ChunkSizes = 43200 ;
		ted_pro_tel0_hi_eflux:_DeflateLevel = 9 ;
		ted_pro_tel0_hi_eflux:_Shuffle = "true" ;
		ted_pro_tel0_hi_eflux:_FillValue = -1e+31 ;
	float ted_pro_tel30_hi_eflux(time) ;
		ted_pro_tel30_hi_eflux:long_name = "TED proton (1-20 keV)  30 deg telescope energy flux" ;
		ted_pro_tel30_hi_eflux:units = "mW/m2-str" ;
		ted_pro_tel30_hi_eflux:valid_range = -200., 200. ;
		ted_pro_tel30_hi_eflux:_Storage = "chunked" ;
		ted_pro_tel30_hi_eflux:_ChunkSizes = 43200 ;
		ted_pro_tel30_hi_eflux:_DeflateLevel = 9 ;
		ted_pro_tel30_hi_eflux:_Shuffle = "true" ;
		ted_pro_tel30_hi_eflux:_FillValue = -1e+31 ;
	int ted_ele_tel0_low_eflux_error(time) ;
		ted_ele_tel0_low_eflux_error:long_name = "TED electron (50eV-1 keV) 0 deg telescope energy flux percent error" ;
		ted_ele_tel0_low_eflux_error:units = "mW/m2-str" ;
		ted_ele_tel0_low_eflux_error:_Storage = "chunked" ;
		ted_ele_tel0_low_eflux_error:_ChunkSizes = 43200 ;
		ted_ele_tel0_low_eflux_error:_DeflateLevel = 9 ;
		ted_ele_tel0_low_eflux_error:_Shuffle = "true" ;
		ted_ele_tel0_low_eflux_error:_Endianness = "little" ;
		ted_ele_tel0_low_eflux_error:_FillValue = -2147483647 ;
	int ted_ele_tel30_low_eflux_error(time) ;
		ted_ele_tel30_low_eflux_error:long_name = "TED electron (50eV-1 keV) 30 deg telescope energy flux percent error" ;
		ted_ele_tel30_low_eflux_error:units = "mW/m2-str" ;
		ted_ele_tel30_low_eflux_error:_Storage = "chunked" ;
		ted_ele_tel30_low_eflux_error:_ChunkSizes = 43200 ;
		ted_ele_tel30_low_eflux_error:_DeflateLevel = 9 ;
		ted_ele_tel30_low_eflux_error:_Shuffle = "true" ;
		ted_ele_tel30_low_eflux_error:_Endianness = "little" ;
		ted_ele_tel30_low_eflux_error:_FillValue = -2147483647 ;
	int ted_ele_tel0_hi_eflux_error(time) ;
		ted_ele_tel0_hi_eflux_error:long_name = "TED electron (1-20 keV) 0 deg telescope energy flux percent error" ;
		ted_ele_tel0_hi_eflux_error:units = "mW/m2-str" ;
		ted_ele_tel0_hi_eflux_error:_Storage = "chunked" ;
		ted_ele_tel0_hi_eflux_error:_ChunkSizes = 43200 ;
		ted_ele_tel0_hi_eflux_error:_DeflateLevel = 9 ;
		ted_ele_tel0_hi_eflux_error:_Shuffle = "true" ;
		ted_ele_tel0_hi_eflux_error:_Endianness = "little" ;
		ted_ele_tel0_hi_eflux_error:_FillValue = -2147483647 ;
	int ted_ele_tel30_hi_eflux_error(time) ;
		ted_ele_tel30_hi_eflux_error:long_name = "TED electron (1-20 keV)  30 deg telescope energy flux percent error" ;
		ted_ele_tel30_hi_eflux_error:units = "mW/m2-str" ;
		ted_ele_tel30_hi_eflux_error:_Storage = "chunked" ;
		ted_ele_tel30_hi_eflux_error:_ChunkSizes = 43200 ;
		ted_ele_tel30_hi_eflux_error:_DeflateLevel = 9 ;
		ted_ele_tel30_hi_eflux_error:_Shuffle = "true" ;
		ted_ele_tel30_hi_eflux_error:_Endianness = "little" ;
		ted_ele_tel30_hi_eflux_error:_FillValue = -2147483647 ;
	int ted_pro_tel0_low_eflux_error(time) ;
		ted_pro_tel0_low_eflux_error:long_name = "TED proton (50eV-1 keV) 0 deg telescope energy flux percent error" ;
		ted_pro_tel0_low_eflux_error:units = "mW/m2-str" ;
		ted_pro_tel0_low_eflux_error:_Storage = "chunked" ;
		ted_pro_tel0_low_eflux_error:_ChunkSizes = 43200 ;
		ted_pro_tel0_low_eflux_error:_DeflateLevel = 9 ;
		ted_pro_tel0_low_eflux_error:_Shuffle = "true" ;
		ted_pro_tel0_low_eflux_error:_Endianness = "little" ;
		ted_pro_tel0_low_eflux_error:_FillValue = -2147483647 ;
	int ted_pro_tel30_low_eflux_error(time) ;
		ted_pro_tel30_low_eflux_error:long_name = "TEDproton (50eV-1 keV) 30 deg telescope energy flux percent error" ;
		ted_pro_tel30_low_eflux_error:units = "mW/m2-str" ;
		ted_pro_tel30_low_eflux_error:_Storage = "chunked" ;
		ted_pro_tel30_low_eflux_error:_ChunkSizes = 43200 ;
		ted_pro_tel30_low_eflux_error:_DeflateLevel = 9 ;
		ted_pro_tel30_low_eflux_error:_Shuffle = "true" ;
		ted_pro_tel30_low_eflux_error:_Endianness = "little" ;
		ted_pro_tel30_low_eflux_error:_FillValue = -2147483647 ;
	int ted_pro_tel0_hi_eflux_error(time) ;
		ted_pro_tel0_hi_eflux_error:long_name = "TED proton (1-20 keV)  0 deg telescope energy flux percent error" ;
		ted_pro_tel0_hi_eflux_error:units = "mW/m2-str" ;
		ted_pro_tel0_hi_eflux_error:_Storage = "chunked" ;
		ted_pro_tel0_hi_eflux_error:_ChunkSizes = 43200 ;
		ted_pro_tel0_hi_eflux_error:_DeflateLevel = 9 ;
		ted_pro_tel0_hi_eflux_error:_Shuffle = "true" ;
		ted_pro_tel0_hi_eflux_error:_Endianness = "little" ;
		ted_pro_tel0_hi_eflux_error:_FillValue = -2147483647 ;
	int ted_pro_tel30_hi_eflux_error(time) ;
		ted_pro_tel30_hi_eflux_error:long_name = "TED proton (1-20 keV)  30 deg telescope energy flux percent error" ;
		ted_pro_tel30_hi_eflux_error:units = "mW/m2-str" ;
		ted_pro_tel30_hi_eflux_error:_Storage = "chunked" ;
		ted_pro_tel30_hi_eflux_error:_ChunkSizes = 43200 ;
		ted_pro_tel30_hi_eflux_error:_DeflateLevel = 9 ;
		ted_pro_tel30_hi_eflux_error:_Shuffle = "true" ;
		ted_pro_tel30_hi_eflux_error:_Endianness = "little" ;
		ted_pro_tel30_hi_eflux_error:_FillValue = -2147483647 ;
	float ted_ele_eflux_atmo_low(time) ;
		ted_ele_eflux_atmo_low:long_name = "TED electron (50eV-1 keV) energy flux at 120 km" ;
		ted_ele_eflux_atmo_low:units = "mW/m2" ;
		ted_ele_eflux_atmo_low:valid_range = -6400., 6400. ;
		ted_ele_eflux_atmo_low:_Storage = "chunked" ;
		ted_ele_eflux_atmo_low:_ChunkSizes = 43200 ;
		ted_ele_eflux_atmo_low:_DeflateLevel = 9 ;
		ted_ele_eflux_atmo_low:_Shuffle = "true" ;
		ted_ele_eflux_atmo_low:_FillValue = -1e+31 ;
	float ted_ele_eflux_atmo_hi(time) ;
		ted_ele_eflux_atmo_hi:long_name = "TED electron (1-20 keV) energy flux at 120 km" ;
		ted_ele_eflux_atmo_hi:units = "mW/m2" ;
		ted_ele_eflux_atmo_hi:valid_range = -6400., 6400. ;
		ted_ele_eflux_atmo_hi:_Storage = "chunked" ;
		ted_ele_eflux_atmo_hi:_ChunkSizes = 43200 ;
		ted_ele_eflux_atmo_hi:_DeflateLevel = 9 ;
		ted_ele_eflux_atmo_hi:_Shuffle = "true" ;
		ted_ele_eflux_atmo_hi:_FillValue = -1e+31 ;
	float ted_ele_eflux_atmo_total(time) ;
		ted_ele_eflux_atmo_total:long_name = "TED electron (50 eV-20 keV) energy flux at 120 km" ;
		ted_ele_eflux_atmo_total:units = "mW/m2" ;
		ted_ele_eflux_atmo_total:valid_range = -12800., 6400. ;
		ted_ele_eflux_atmo_total:_Storage = "chunked" ;
		ted_ele_eflux_atmo_total:_ChunkSizes = 43200 ;
		ted_ele_eflux_atmo_total:_DeflateLevel = 9 ;
		ted_ele_eflux_atmo_total:_Shuffle = "true" ;
		ted_ele_eflux_atmo_total:_FillValue = -1e+31 ;
	int ted_ele_eflux_atmo_low_err(time) ;
		ted_ele_eflux_atmo_low_err:long_name = "TED electron (50eV-1 keV) energy flux percent error at 120 km" ;
		ted_ele_eflux_atmo_low_err:units = "mW/m2" ;
		ted_ele_eflux_atmo_low_err:valid_range = 0., 6400. ;
		ted_ele_eflux_atmo_low_err:_Storage = "chunked" ;
		ted_ele_eflux_atmo_low_err:_ChunkSizes = 43200 ;
		ted_ele_eflux_atmo_low_err:_DeflateLevel = 9 ;
		ted_ele_eflux_atmo_low_err:_Shuffle = "true" ;
		ted_ele_eflux_atmo_low_err:_Endianness = "little" ;
		ted_ele_eflux_atmo_low_err:_FillValue = -2147483647 ;
	int ted_ele_eflux_atmo_hi_err(time) ;
		ted_ele_eflux_atmo_hi_err:long_name = "TED electron (1-20 keV) energy flux percent error at 120 km" ;
		ted_ele_eflux_atmo_hi_err:units = "mW/m2" ;
		ted_ele_eflux_atmo_hi_err:valid_range = 0., 6400. ;
		ted_ele_eflux_atmo_hi_err:_Storage = "chunked" ;
		ted_ele_eflux_atmo_hi_err:_ChunkSizes = 43200 ;
		ted_ele_eflux_atmo_hi_err:_DeflateLevel = 9 ;
		ted_ele_eflux_atmo_hi_err:_Shuffle = "true" ;
		ted_ele_eflux_atmo_hi_err:_Endianness = "little" ;
		ted_ele_eflux_atmo_hi_err:_FillValue = -2147483647 ;
	int ted_ele_eflux_atmo_total_err(time) ;
		ted_ele_eflux_atmo_total_err:long_name = "TED electron (50 eV-20 keV) energy flux percent error at 120 km" ;
		ted_ele_eflux_atmo_total_err:units = "mW/m2" ;
		ted_ele_eflux_atmo_total_err:valid_range = 0., 6400. ;
		ted_ele_eflux_atmo_total_err:_Storage = "chunked" ;
		ted_ele_eflux_atmo_total_err:_ChunkSizes = 43200 ;
		ted_ele_eflux_atmo_total_err:_DeflateLevel = 9 ;
		ted_ele_eflux_atmo_total_err:_Shuffle = "true" ;
		ted_ele_eflux_atmo_total_err:_Endianness = "little" ;
		ted_ele_eflux_atmo_total_err:_FillValue = -2147483647 ;
	float ted_pro_eflux_atmo_low(time) ;
		ted_pro_eflux_atmo_low:long_name = "TED proton (50eV-1 keV) energy flux at 120 km" ;
		ted_pro_eflux_atmo_low:units = "mW/m2" ;
		ted_pro_eflux_atmo_low:valid_range = -6400., 6400. ;
		ted_pro_eflux_atmo_low:_Storage = "chunked" ;
		ted_pro_eflux_atmo_low:_ChunkSizes = 43200 ;
		ted_pro_eflux_atmo_low:_DeflateLevel = 9 ;
		ted_pro_eflux_atmo_low:_Shuffle = "true" ;
		ted_pro_eflux_atmo_low:_FillValue = -1e+31 ;
	float ted_pro_eflux_atmo_hi(time) ;
		ted_pro_eflux_atmo_hi:long_name = "TED proton (1-20 keV) energy flux at 120 km" ;
		ted_pro_eflux_atmo_hi:units = "mW/m2" ;
		ted_pro_eflux_atmo_hi:valid_range = -6400., 6400. ;
		ted_pro_eflux_atmo_hi:_Storage = "chunked" ;
		ted_pro_eflux_atmo_hi:_ChunkSizes = 43200 ;
		ted_pro_eflux_atmo_hi:_DeflateLevel = 9 ;
		ted_pro_eflux_atmo_hi:_Shuffle = "true" ;
		ted_pro_eflux_atmo_hi:_FillValue = -1e+31 ;
	float ted_pro_eflux_atmo_total(time) ;
		ted_pro_eflux_atmo_total:long_name = "TED proton (50 eV-20 keV) energy flux at 120 km" ;
		ted_pro_eflux_atmo_total:units = "mW/m2" ;
		ted_pro_eflux_atmo_total:valid_range = -12800., 12800. ;
		ted_pro_eflux_atmo_total:_Storage = "chunked" ;
		ted_pro_eflux_atmo_total:_ChunkSizes = 43200 ;
		ted_pro_eflux_atmo_total:_DeflateLevel = 9 ;
		ted_pro_eflux_atmo_total:_Shuffle = "true" ;
		ted_pro_eflux_atmo_total:_FillValue = -1e+31 ;
	int ted_pro_eflux_atmo_low_err(time) ;
		ted_pro_eflux_atmo_low_err:long_name = "TED proton (50eV-1 keV) energy flux percent error at 120 km" ;
		ted_pro_eflux_atmo_low_err:units = "mW/m2" ;
		ted_pro_eflux_atmo_low_err:valid_range = 0., 6400. ;
		ted_pro_eflux_atmo_low_err:_Storage = "chunked" ;
		ted_pro_eflux_atmo_low_err:_ChunkSizes = 43200 ;
		ted_pro_eflux_atmo_low_err:_DeflateLevel = 9 ;
		ted_pro_eflux_atmo_low_err:_Shuffle = "true" ;
		ted_pro_eflux_atmo_low_err:_Endianness = "little" ;
		ted_pro_eflux_atmo_low_err:_FillValue = -2147483647 ;
	int ted_pro_eflux_atmo_hi_err(time) ;
		ted_pro_eflux_atmo_hi_err:long_name = "TED proton (1-20 keV) energy flux percent error at 120 km" ;
		ted_pro_eflux_atmo_hi_err:units = "mW/m2" ;
		ted_pro_eflux_atmo_hi_err:valid_range = 0., 6400. ;
		ted_pro_eflux_atmo_hi_err:_Storage = "chunked" ;
		ted_pro_eflux_atmo_hi_err:_ChunkSizes = 43200 ;
		ted_pro_eflux_atmo_hi_err:_DeflateLevel = 9 ;
		ted_pro_eflux_atmo_hi_err:_Shuffle = "true" ;
		ted_pro_eflux_atmo_hi_err:_Endianness = "little" ;
		ted_pro_eflux_atmo_hi_err:_FillValue = -2147483647 ;
	int ted_pro_eflux_atmo_total_err(time) ;
		ted_pro_eflux_atmo_total_err:long_name = "TED proton (50 eV-20 keV) energy flux percent error at 120 km" ;
		ted_pro_eflux_atmo_total_err:units = "mW/m2" ;
		ted_pro_eflux_atmo_total_err:valid_range = 0., 12800. ;
		ted_pro_eflux_atmo_total_err:_Storage = "chunked" ;
		ted_pro_eflux_atmo_total_err:_ChunkSizes = 43200 ;
		ted_pro_eflux_atmo_total_err:_DeflateLevel = 9 ;
		ted_pro_eflux_atmo_total_err:_Shuffle = "true" ;
		ted_pro_eflux_atmo_total_err:_Endianness = "little" ;
		ted_pro_eflux_atmo_total_err:_FillValue = -2147483647 ;
	float ted_total_eflux_atmo(time) ;
		ted_total_eflux_atmo:long_name = "TED total (50 ev-20 keV) energy flux of protons and electrons at 120 km" ;
		ted_total_eflux_atmo:units = "mW/m2" ;
		ted_total_eflux_atmo:valid_range = -25600., 25600. ;
		ted_total_eflux_atmo:_Storage = "chunked" ;
		ted_total_eflux_atmo:_ChunkSizes = 43200 ;
		ted_total_eflux_atmo:_DeflateLevel = 9 ;
		ted_total_eflux_atmo:_Shuffle = "true" ;
		ted_total_eflux_atmo:_FillValue = -1e+31 ;
	int ted_total_eflux_atmo_err(time) ;
		ted_total_eflux_atmo_err:long_name = "TED total (50 ev-20 keV) energy flux percent error of protons and electrons at 120 km" ;
		ted_total_eflux_atmo_err:units = "mW/m2" ;
		ted_total_eflux_atmo_err:valid_range = -25600., 25600. ;
		ted_total_eflux_atmo_err:_Storage = "chunked" ;
		ted_total_eflux_atmo_err:_ChunkSizes = 43200 ;
		ted_total_eflux_atmo_err:_DeflateLevel = 9 ;
		ted_total_eflux_atmo_err:_Shuffle = "true" ;
		ted_total_eflux_atmo_err:_Endianness = "little" ;
		ted_total_eflux_atmo_err:_FillValue = -2147483647 ;
	byte ted_ele_energy_tel0(time) ;
		ted_ele_energy_tel0:long_name = "TED electron characteristic energy channel 0 deg telescope" ;
		ted_ele_energy_tel0:units = "energy channel" ;
		ted_ele_energy_tel0:valid_range = 0., 15. ;
		ted_ele_energy_tel0:_Storage = "chunked" ;
		ted_ele_energy_tel0:_ChunkSizes = 43200 ;
		ted_ele_energy_tel0:_DeflateLevel = 9 ;
		ted_ele_energy_tel0:_Shuffle = "true" ;
	byte ted_ele_energy_tel30(time) ;
		ted_ele_energy_tel30:long_name = "TED electron characteristic energy channel 30 deg telescope" ;
		ted_ele_energy_tel30:units = "energy channel" ;
		ted_ele_energy_tel30:valid_range = 0., 15. ;
		ted_ele_energy_tel30:_Storage = "chunked" ;
		ted_ele_energy_tel30:_ChunkSizes = 43200 ;
		ted_ele_energy_tel30:_DeflateLevel = 9 ;
		ted_ele_energy_tel30:_Shuffle = "true" ;
	byte ted_pro_energy_tel0(time) ;
		ted_pro_energy_tel0:long_name = "TED proton characteristic energy channel  0 deg telescope" ;
		ted_pro_energy_tel0:units = "energy channel" ;
		ted_pro_energy_tel0:valid_range = 0., 15. ;
		ted_pro_energy_tel0:_Storage = "chunked" ;
		ted_pro_energy_tel0:_ChunkSizes = 43200 ;
		ted_pro_energy_tel0:_DeflateLevel = 9 ;
		ted_pro_energy_tel0:_Shuffle = "true" ;
	byte ted_pro_energy_tel30(time) ;
		ted_pro_energy_tel30:long_name = "TED proton characteristic energy channel 30 deg telescope" ;
		ted_pro_energy_tel30:units = "energy channel" ;
		ted_pro_energy_tel30:valid_range = 0., 15. ;
		ted_pro_energy_tel30:_Storage = "chunked" ;
		ted_pro_energy_tel30:_ChunkSizes = 43200 ;
		ted_pro_energy_tel30:_DeflateLevel = 9 ;
		ted_pro_energy_tel30:_Shuffle = "true" ;
	float ted_ele_max_flux_tel0(time) ;
		ted_ele_max_flux_tel0:long_name = "TED electron maximum flux [#/cm2-s-str-eV] 0 deg telescope" ;
		ted_ele_max_flux_tel0:units = "[#/cm2-s-str-eV]" ;
		ted_ele_max_flux_tel0:valid_range = 0., 4000000000. ;
		ted_ele_max_flux_tel0:_Storage = "chunked" ;
		ted_ele_max_flux_tel0:_ChunkSizes = 43200 ;
		ted_ele_max_flux_tel0:_DeflateLevel = 9 ;
		ted_ele_max_flux_tel0:_Shuffle = "true" ;
		ted_ele_max_flux_tel0:_FillValue = -1e+31 ;
	float ted_ele_max_flux_tel30(time) ;
		ted_ele_max_flux_tel30:long_name = "TED electron maximum flux [#/cm2-s-str-eV] 30 deg telescope" ;
		ted_ele_max_flux_tel30:units = "[#/cm2-s-str-eV]" ;
		ted_ele_max_flux_tel30:valid_range = 0., 4000000000. ;
		ted_ele_max_flux_tel30:_Storage = "chunked" ;
		ted_ele_max_flux_tel30:_ChunkSizes = 43200 ;
		ted_ele_max_flux_tel30:_DeflateLevel = 9 ;
		ted_ele_max_flux_tel30:_Shuffle = "true" ;
		ted_ele_max_flux_tel30:_FillValue = -1e+31 ;
	float ted_pro_max_flux_tel0(time) ;
		ted_pro_max_flux_tel0:long_name = "TED proton maximum flux [#/cm2-s-str-eV] 0 deg telescope" ;
		ted_pro_max_flux_tel0:units = "[#/cm2-s-str-eV" ;
		ted_pro_max_flux_tel0:valid_range = 0., 4000000000. ;
		ted_pro_max_flux_tel0:_Storage = "chunked" ;
		ted_pro_max_flux_tel0:_ChunkSizes = 43200 ;
		ted_pro_max_flux_tel0:_DeflateLevel = 9 ;
		ted_pro_max_flux_tel0:_Shuffle = "true" ;
		ted_pro_max_flux_tel0:_FillValue = -1e+31 ;
	float ted_pro_max_flux_tel30(time) ;
		ted_pro_max_flux_tel30:long_name = "TED proton maximum flux [#/cm2-s-str-eV] 30 deg telescope" ;
		ted_pro_max_flux_tel30:units = "[#/cm2-s-str-eV" ;
		ted_pro_max_flux_tel30:valid_range = 0., 4000000000. ;
		ted_pro_max_flux_tel30:_Storage = "chunked" ;
		ted_pro_max_flux_tel30:_ChunkSizes = 43200 ;
		ted_pro_max_flux_tel30:_DeflateLevel = 9 ;
		ted_pro_max_flux_tel30:_Shuffle = "true" ;
		ted_pro_max_flux_tel30:_FillValue = -1e+31 ;
	float ted_ele_eflux_bg_tel0_low(time) ;
		ted_ele_eflux_bg_tel0_low:long_name = "TED electron background low energy 0 degree telescope" ;
		ted_ele_eflux_bg_tel0_low:units = "mW/m2-str" ;
		ted_ele_eflux_bg_tel0_low:valid_range = 0., 200. ;
		ted_ele_eflux_bg_tel0_low:_Storage = "chunked" ;
		ted_ele_eflux_bg_tel0_low:_ChunkSizes = 43200 ;
		ted_ele_eflux_bg_tel0_low:_DeflateLevel = 9 ;
		ted_ele_eflux_bg_tel0_low:_Shuffle = "true" ;
		ted_ele_eflux_bg_tel0_low:_FillValue = -1e+31 ;
	float ted_ele_eflux_bg_tel30_low(time) ;
		ted_ele_eflux_bg_tel30_low:long_name = "TED electron background low energy 30 degree telescope" ;
		ted_ele_eflux_bg_tel30_low:units = "mW/m2-str" ;
		ted_ele_eflux_bg_tel30_low:valid_range = 0., 200. ;
		ted_ele_eflux_bg_tel30_low:_Storage = "chunked" ;
		ted_ele_eflux_bg_tel30_low:_ChunkSizes = 43200 ;
		ted_ele_eflux_bg_tel30_low:_DeflateLevel = 9 ;
		ted_ele_eflux_bg_tel30_low:_Shuffle = "true" ;
		ted_ele_eflux_bg_tel30_low:_FillValue = -1e+31 ;
	float ted_ele_eflux_bg_tel0_hi(time) ;
		ted_ele_eflux_bg_tel0_hi:long_name = "TED electron background high energy 0 degree telescope" ;
		ted_ele_eflux_bg_tel0_hi:units = "mW/m2-str" ;
		ted_ele_eflux_bg_tel0_hi:valid_range = 0., 200. ;
		ted_ele_eflux_bg_tel0_hi:_Storage = "chunked" ;
		ted_ele_eflux_bg_tel0_hi:_ChunkSizes = 43200 ;
		ted_ele_eflux_bg_tel0_hi:_DeflateLevel = 9 ;
		ted_ele_eflux_bg_tel0_hi:_Shuffle = "true" ;
		ted_ele_eflux_bg_tel0_hi:_FillValue = -1e+31 ;
	float ted_ele_eflux_bg_tel30_hi(time) ;
		ted_ele_eflux_bg_tel30_hi:long_name = "TED electron background high energy 30 degree telescope" ;
		ted_ele_eflux_bg_tel30_hi:units = "mW/m2-str" ;
		ted_ele_eflux_bg_tel30_hi:valid_range = 0., 200. ;
		ted_ele_eflux_bg_tel30_hi:_Storage = "chunked" ;
		ted_ele_eflux_bg_tel30_hi:_ChunkSizes = 43200 ;
		ted_ele_eflux_bg_tel30_hi:_DeflateLevel = 9 ;
		ted_ele_eflux_bg_tel30_hi:_Shuffle = "true" ;
		ted_ele_eflux_bg_tel30_hi:_FillValue = -1e+31 ;
	float ted_pro_eflux_bg_tel0_low(time) ;
		ted_pro_eflux_bg_tel0_low:long_name = "TED proton background low energy 0 degree telescope" ;
		ted_pro_eflux_bg_tel0_low:units = "mW/m2-str" ;
		ted_pro_eflux_bg_tel0_low:valid_range = 0., 200. ;
		ted_pro_eflux_bg_tel0_low:_Storage = "chunked" ;
		ted_pro_eflux_bg_tel0_low:_ChunkSizes = 43200 ;
		ted_pro_eflux_bg_tel0_low:_DeflateLevel = 9 ;
		ted_pro_eflux_bg_tel0_low:_Shuffle = "true" ;
		ted_ele_eflux_bg_tel0_low:_FillValue = -1e+31 ;
	float ted_pro_eflux_bg_tel30_low(time) ;
		ted_pro_eflux_bg_tel30_low:long_name = "TED proton background low energy 30 degree telescope" ;
		ted_pro_eflux_bg_tel30_low:units = "mW/m2-str" ;
		ted_pro_eflux_bg_tel30_low:valid_range = 0., 200. ;
		ted_pro_eflux_bg_tel30_low:_Storage = "chunked" ;
		ted_pro_eflux_bg_tel30_low:_ChunkSizes = 43200 ;
		ted_pro_eflux_bg_tel30_low:_DeflateLevel = 9 ;
		ted_pro_eflux_bg_tel30_low:_Shuffle = "true" ;
		ted_ele_eflux_bg_tel30_low:_FillValue = -1e+31 ;
	float ted_pro_eflux_bg_tel0_hi(time) ;
		ted_pro_eflux_bg_tel0_hi:long_name = "TED proton background high energy 0 degree telescope" ;
		ted_pro_eflux_bg_tel0_hi:units = "mW/m2-str" ;
		ted_pro_eflux_bg_tel0_hi:valid_range = 0., 200. ;
		ted_pro_eflux_bg_tel0_hi:_Storage = "chunked" ;
		ted_pro_eflux_bg_tel0_hi:_ChunkSizes = 43200 ;
		ted_pro_eflux_bg_tel0_hi:_DeflateLevel = 9 ;
		ted_pro_eflux_bg_tel0_hi:_Shuffle = "true" ;
		ted_ele_eflux_bg_tel0_hi:_FillValue = -1e+31 ;
	float ted_pro_eflux_bg_tel30_hi(time) ;
		ted_pro_eflux_bg_tel30_hi:long_name = "TED proton background high energy 30 degree telescope" ;
		ted_pro_eflux_bg_tel30_hi:units = "mW/m2-str" ;
		ted_pro_eflux_bg_tel30_hi:valid_range = 0., 200. ;
		ted_pro_eflux_bg_tel30_hi:_Storage = "chunked" ;
		ted_pro_eflux_bg_tel30_hi:_ChunkSizes = 43200 ;
		ted_pro_eflux_bg_tel30_hi:_DeflateLevel = 9 ;
		ted_pro_eflux_bg_tel30_hi:_Shuffle = "true" ;
		ted_ele_eflux_bg_tel30_hi:_FillValue = -1e+31 ;
	float ted_ele_eflux_bg_tel0_low_cps(time) ;
		ted_ele_eflux_bg_tel0_low_cps:long_name = "TED electron background low energy 0 degree telescope counts" ;
		ted_ele_eflux_bg_tel0_low_cps:units = "counts" ;
		ted_ele_eflux_bg_tel0_low_cps:valid_range = 0., 1998848. ;
		ted_ele_eflux_bg_tel0_low_cps:_Storage = "chunked" ;
		ted_ele_eflux_bg_tel0_low_cps:_ChunkSizes = 43200 ;
		ted_ele_eflux_bg_tel0_low_cps:_DeflateLevel = 9 ;
		ted_ele_eflux_bg_tel0_low_cps:_Shuffle = "true" ;
		ted_ele_eflux_bg_tel0_low:_FillValue = -1e+31 ;
	float ted_ele_eflux_bg_tel30_low_cps(time) ;
		ted_ele_eflux_bg_tel30_low_cps:long_name = "TED electron background low energy 30 degree telescope counts" ;
		ted_ele_eflux_bg_tel30_low_cps:units = "counts" ;
		ted_ele_eflux_bg_tel30_low_cps:valid_range = 0., 1998848. ;
		ted_ele_eflux_bg_tel30_low_cps:_Storage = "chunked" ;
		ted_ele_eflux_bg_tel30_low_cps:_ChunkSizes = 43200 ;
		ted_ele_eflux_bg_tel30_low_cps:_DeflateLevel = 9 ;
		ted_ele_eflux_bg_tel30_low_cps:_Shuffle = "true" ;
		ted_ele_eflux_bg_tel30_low:_FillValue = -1e+31 ;
	float ted_ele_eflux_bg_tel0_hi_cps(time) ;
		ted_ele_eflux_bg_tel0_hi_cps:long_name = "TED electron background high energy 0 degree telescope counts" ;
		ted_ele_eflux_bg_tel0_hi_cps:units = "counts" ;
		ted_ele_eflux_bg_tel0_hi_cps:valid_range = 0., 1998848. ;
		ted_ele_eflux_bg_tel0_hi_cps:_Storage = "chunked" ;
		ted_ele_eflux_bg_tel0_hi_cps:_ChunkSizes = 43200 ;
		ted_ele_eflux_bg_tel0_hi_cps:_DeflateLevel = 9 ;
		ted_ele_eflux_bg_tel0_hi_cps:_Shuffle = "true" ;
		ted_ele_eflux_bg_tel0_hi:_FillValue = -1e+31 ;
	float ted_ele_eflux_bg_tel30_hi_cps(time) ;
		ted_ele_eflux_bg_tel30_hi_cps:long_name = "TED electron background high energy 30 degree telescope counts" ;
		ted_ele_eflux_bg_tel30_hi_cps:units = "counts" ;
		ted_ele_eflux_bg_tel30_hi_cps:valid_range = 0., 1998848. ;
		ted_ele_eflux_bg_tel30_hi_cps:_Storage = "chunked" ;
		ted_ele_eflux_bg_tel30_hi_cps:_ChunkSizes = 43200 ;
		ted_ele_eflux_bg_tel30_hi_cps:_DeflateLevel = 9 ;
		ted_ele_eflux_bg_tel30_hi_cps:_Shuffle = "true" ;
		ted_ele_eflux_bg_tel30_hi:_FillValue = -1e+31 ;
	float ted_pro_eflux_bg_tel0_low_cps(time) ;
		ted_pro_eflux_bg_tel0_low_cps:long_name = "TED proton background low energy 0 degree telescope counts" ;
		ted_pro_eflux_bg_tel0_low_cps:units = "counts" ;
		ted_pro_eflux_bg_tel0_low_cps:valid_range = 0., 1998848. ;
		ted_pro_eflux_bg_tel0_low_cps:_Storage = "chunked" ;
		ted_pro_eflux_bg_tel0_low_cps:_ChunkSizes = 43200 ;
		ted_pro_eflux_bg_tel0_low_cps:_DeflateLevel = 9 ;
		ted_pro_eflux_bg_tel0_low_cps:_Shuffle = "true" ;
		ted_pro_eflux_bg_tel0_low_cps:_FillValue = -1e+31 ;
	float ted_pro_eflux_bg_tel30_low_cps(time) ;
		ted_pro_eflux_bg_tel30_low_cps:long_name = "TED proton background low energy 30 degree telescope counts" ;
		ted_pro_eflux_bg_tel30_low_cps:units = "counts" ;
		ted_pro_eflux_bg_tel30_low_cps:valid_range = 0., 1998848. ;
		ted_pro_eflux_bg_tel30_low_cps:_Storage = "chunked" ;
		ted_pro_eflux_bg_tel30_low_cps:_ChunkSizes = 43200 ;
		ted_pro_eflux_bg_tel30_low_cps:_DeflateLevel = 9 ;
		ted_pro_eflux_bg_tel30_low_cps:_Shuffle = "true" ;
		ted_pro_eflux_bg_tel30_low_cps:_FillValue = -1e+31 ;
	float ted_pro_eflux_bg_tel0_hi_cps(time) ;
		ted_pro_eflux_bg_tel0_hi_cps:long_name = "TED proton background high energy 0 degree telescope counts" ;
		ted_pro_eflux_bg_tel0_hi_cps:units = "counts" ;
		ted_pro_eflux_bg_tel0_hi_cps:valid_range = 0., 1998848. ;
		ted_pro_eflux_bg_tel0_hi_cps:_Storage = "chunked" ;
		ted_pro_eflux_bg_tel0_hi_cps:_ChunkSizes = 43200 ;
		ted_pro_eflux_bg_tel0_hi_cps:_DeflateLevel = 9 ;
		ted_pro_eflux_bg_tel0_hi_cps:_Shuffle = "true" ;
		ted_pro_eflux_bg_tel0_hi_cps:_FillValue = -1e+31 ;
	float ted_pro_eflux_bg_tel30_hi_cps(time) ;
		ted_pro_eflux_bg_tel30_hi_cps:long_name = "TED proton background high energy 30 degree telescope counts" ;
		ted_pro_eflux_bg_tel30_hi_cps:units = "counts" ;
		ted_pro_eflux_bg_tel30_hi_cps:valid_range = 0., 1998848. ;
		ted_pro_eflux_bg_tel30_hi_cps:_Storage = "chunked" ;
		ted_pro_eflux_bg_tel30_hi_cps:_ChunkSizes = 43200 ;
		ted_pro_eflux_bg_tel30_hi_cps:_DeflateLevel = 9 ;
		ted_pro_eflux_bg_tel30_hi_cps:_Shuffle = "true" ;
		ted_pro_eflux_bg_tel30_hi_cps:_FillValue = -1e+31 ;
	float Br_sat(time) ;
		Br_sat:long_name = "Bradial IGRF (satellite)" ;
		Br_sat:units = "nT" ;
		Br_sat:valid_range = -50000., 50000. ;
		Br_sat:_Storage = "chunked" ;
		Br_sat:_ChunkSizes = 43200 ;
		Br_sat:_DeflateLevel = 9 ;
		Br_sat:_Shuffle = "true" ;
		Br_sat:_FillValue = -1e+31 ;
	float Bt_sat(time) ;
		Bt_sat:long_name = "Btheta IGRF (satellite)" ;
		Bt_sat:units = "nT" ;
		Bt_sat:valid_range = -50000., 50000. ;
		Bt_sat:_Storage = "chunked" ;
		Bt_sat:_ChunkSizes = 43200 ;
		Bt_sat:_DeflateLevel = 9 ;
		Bt_sat:_Shuffle = "true" ;
		Bt_sat:_FillValue = -1e+31 ;
	float Bp_sat(time) ;
		Bp_sat:long_name = "Bphi IGRF (satellite)" ;
		Bp_sat:units = "nT" ;
		Bp_sat:valid_range = -50000., 50000. ;
		Bp_sat:_Storage = "chunked" ;
		Bp_sat:_ChunkSizes = 43200 ;
		Bp_sat:_DeflateLevel = 9 ;
		Bp_sat:_Shuffle = "true" ;
		Bp_sat:_FillValue = -1e+31 ;
	float Btot_sat(time) ;
		Btot_sat:long_name = "Btotal IGRF (satellite)" ;
		Btot_sat:units = "nT" ;
		Btot_sat:valid_range = -50000., 50000. ;
		Btot_sat:_Storage = "chunked" ;
		Btot_sat:_ChunkSizes = 43200 ;
		Btot_sat:_DeflateLevel = 9 ;
		Btot_sat:_Shuffle = "true" ;
		Btot_sat:_FillValue = -1e+31 ;
	float Br_foot(time) ;
		Br_foot:long_name = "Bradial IGRF (foot of field line)" ;
		Br_foot:units = "nT" ;
		Br_foot:valid_range = -50000., 50000. ;
		Br_foot:_Storage = "chunked" ;
		Br_foot:_ChunkSizes = 43200 ;
		Br_foot:_DeflateLevel = 9 ;
		Br_foot:_Shuffle = "true" ;
		Br_foot:_FillValue = -1e+31 ;
	float Bt_foot(time) ;
		Bt_foot:long_name = "Btheta IGRF (foot of field line)" ;
		Bt_foot:units = "nT" ;
		Bt_foot:valid_range = -50000., 50000. ;
		Bt_foot:_Storage = "chunked" ;
		Bt_foot:_ChunkSizes = 43200 ;
		Bt_foot:_DeflateLevel = 9 ;
		Bt_foot:_Shuffle = "true" ;
		Bt_foot:_FillValue = -1e+31 ;
	float Bp_foot(time) ;
		Bp_foot:long_name = "Bphi IGRF (foot of field line)" ;
		Bp_foot:units = "nT" ;
		Bp_foot:valid_range = -50000., 50000. ;
		Bp_foot:_Storage = "chunked" ;
		Bp_foot:_ChunkSizes = 43200 ;
		Bp_foot:_DeflateLevel = 9 ;
		Bp_foot:_Shuffle = "true" ;
		Bp_foot:_FillValue = -1e+31 ;
	float Btot_foot(time) ;
		Btot_foot:long_name = "Btotal IGRF (foot of field line)" ;
		Btot_foot:units = "nT" ;
		Btot_foot:valid_range = -50000., 50000. ;
		Btot_foot:_Storage = "chunked" ;
		Btot_foot:_ChunkSizes = 43200 ;
		Btot_foot:_DeflateLevel = 9 ;
		Btot_foot:_Shuffle = "true" ;
		Btot_foot:_FillValue = -1e+31 ;
	float geod_lat_foot(time) ;
		geod_lat_foot:long_name = "Geodetic latitude (foot of field line)" ;
		geod_lat_foot:units = "deg" ;
		geod_lat_foot:valid_range = -90., 90. ;
		geod_lat_foot:_Storage = "chunked" ;
		geod_lat_foot:_ChunkSizes = 43200 ;
		geod_lat_foot:_DeflateLevel = 9 ;
		geod_lat_foot:_Shuffle = "true" ;
		geod_lat_foot:_FillValue = -1e+31 ;
	float geod_lon_foot(time) ;
		geod_lon_foot:long_name = "Geodetic longitude (foot of field line)" ;
		geod_lon_foot:units = "deg" ;
		geod_lon_foot:valid_range = 0., 360. ;
		geod_lon_foot:_Storage = "chunked" ;
		geod_lon_foot:_ChunkSizes = 43200 ;
		geod_lon_foot:_DeflateLevel = 9 ;
		geod_lon_foot:_Shuffle = "true" ;
		geod_lon_foot:_FillValue = -1e+31 ;
	float aacgm_lat_foot(time) ;
		aacgm_lat_foot:long_name = "AACGM latitude (foot of field line)" ;
		aacgm_lat_foot:units = "deg" ;
		aacgm_lat_foot:valid_range = -90., 90. ;
		aacgm_lat_foot:_Storage = "chunked" ;
		aacgm_lat_foot:_ChunkSizes = 43200 ;
		aacgm_lat_foot:_DeflateLevel = 9 ;
		aacgm_lat_foot:_Shuffle = "true" ;
		aacgm_lat_foot:_FillValue = -1e+31 ;
	float aacgm_lon_foot(time) ;
		aacgm_lon_foot:long_name = "AACGM longitude (foot of field line)" ;
		aacgm_lon_foot:units = "deg" ;
		aacgm_lon_foot:valid_range = 0., 360. ;
		aacgm_lon_foot:_Storage = "chunked" ;
		aacgm_lon_foot:_ChunkSizes = 43200 ;
		aacgm_lon_foot:_DeflateLevel = 9 ;
		aacgm_lon_foot:_Shuffle = "true" ;
		aacgm_lon_foot:_FillValue = -1e+31 ;
	float mag_lat_foot(time) ;
		mag_lat_foot:long_name = "magnetic latitude (foot of field line)" ;
		mag_lat_foot:units = "deg" ;
		mag_lat_foot:valid_range = -90., 90. ;
		mag_lat_foot:_Storage = "chunked" ;
		mag_lat_foot:_ChunkSizes = 43200 ;
		mag_lat_foot:_DeflateLevel = 9 ;
		mag_lat_foot:_Shuffle = "true" ;
		mag_lat_foot:_FillValue = -1e+31 ;
	float mag_lon_foot(time) ;
		mag_lon_foot:long_name = "magnetic longitude (foot of field line)" ;
		mag_lon_foot:units = "deg" ;
		mag_lon_foot:valid_range = 0., 360. ;
		mag_lon_foot:_Storage = "chunked" ;
		mag_lon_foot:_ChunkSizes = 43200 ;
		mag_lon_foot:_DeflateLevel = 9 ;
		mag_lon_foot:_Shuffle = "true" ;
		mag_lon_foot:_FillValue = -1e+31 ;
	float mag_lat_sat(time) ;
		mag_lat_sat:long_name = "magnetic latitude (satellite)" ;
		mag_lat_sat:units = "deg" ;
		mag_lat_sat:valid_range = -90., 90. ;
		mag_lat_sat:_Storage = "chunked" ;
		mag_lat_sat:_ChunkSizes = 43200 ;
		mag_lat_sat:_DeflateLevel = 9 ;
		mag_lat_sat:_Shuffle = "true" ;
		mag_lat_sat:_FillValue = -1e+31 ;
	float mag_lon_sat(time) ;
		mag_lon_sat:long_name = "magnetic longitude (satellite)" ;
		mag_lon_sat:units = "deg" ;
		mag_lon_sat:valid_range = 0., 360. ;
		mag_lon_sat:_Storage = "chunked" ;
		mag_lon_sat:_ChunkSizes = 43200 ;
		mag_lon_sat:_DeflateLevel = 9 ;
		mag_lon_sat:_Shuffle = "true" ;
		mag_lon_sat:_FillValue = -1e+31 ;
	float Bx_sat(time) ;
		Bx_sat:long_name = "Bx IGRF satellite coordinates (towards Earth)" ;
		Bx_sat:units = "nT" ;
		Bx_sat:valid_range = -50000., 50000. ;
		Bx_sat:_Storage = "chunked" ;
		Bx_sat:_ChunkSizes = 43200 ;
		Bx_sat:_DeflateLevel = 9 ;
		Bx_sat:_Shuffle = "true" ;
		Bx_sat:_FillValue = -1e+31 ;
	float By_sat(time) ;
		By_sat:long_name = "By IGRF satellite coordinates (opposite velocity direction)" ;
		By_sat:units = "nT" ;
		By_sat:valid_range = -50000., 50000. ;
		By_sat:_Storage = "chunked" ;
		By_sat:_ChunkSizes = 43200 ;
		By_sat:_DeflateLevel = 9 ;
		By_sat:_Shuffle = "true" ;
		By_sat:_FillValue = -1e+31 ;
	float Bz_sat(time) ;
		Bz_sat:long_name = "Bz IGRF satellite coordinates (XxY direction)" ;
		Bz_sat:units = "nT" ;
		Bz_sat:valid_range = -50000., 50000. ;
		Bz_sat:_Storage = "chunked" ;
		Bz_sat:_ChunkSizes = 43200 ;
		Bz_sat:_DeflateLevel = 9 ;
		Bz_sat:_Shuffle = "true" ;
		Bz_sat:_FillValue = -1e+31 ;
	float ted_alpha_0_sat(time) ;
		ted_alpha_0_sat:long_name = "TED 0 deg telescope pitch angle (satellite)" ;
		ted_alpha_0_sat:units = "deg" ;
		ted_alpha_0_sat:valid_range = 0., 180. ;
		ted_alpha_0_sat:_Storage = "chunked" ;
		ted_alpha_0_sat:_ChunkSizes = 43200 ;
		ted_alpha_0_sat:_DeflateLevel = 9 ;
		ted_alpha_0_sat:_Shuffle = "true" ;
		ted_alpha_0_sat:_FillValue = -1e+31 ;
	float ted_alpha_30_sat(time) ;
		ted_alpha_30_sat:long_name = "TED 30 deg telescope pitch angle (satellite)" ;
		ted_alpha_30_sat:units = "deg" ;
		ted_alpha_30_sat:valid_range = 0., 180. ;
		ted_alpha_30_sat:_Storage = "chunked" ;
		ted_alpha_30_sat:_ChunkSizes = 43200 ;
		ted_alpha_30_sat:_DeflateLevel = 9 ;
		ted_alpha_30_sat:_Shuffle = "true" ;
		ted_alpha_30_sat:_FillValue = -1e+31 ;
	float ted_alpha_0_foot(time) ;
		ted_alpha_0_foot:long_name = "TED 0 deg telescope pitch angle (foot of field line)" ;
		ted_alpha_0_foot:units = "deg" ;
		ted_alpha_0_foot:valid_range = 0., 180. ;
		ted_alpha_0_foot:_Storage = "chunked" ;
		ted_alpha_0_foot:_ChunkSizes = 43200 ;
		ted_alpha_0_foot:_DeflateLevel = 9 ;
		ted_alpha_0_foot:_Shuffle = "true" ;
		ted_alpha_0_foot:_FillValue = -1e+31 ;
	float ted_alpha_30_foot(time) ;
		ted_alpha_30_foot:long_name = "TED 30 deg telescope pitch angle (foot of field line)" ;
		ted_alpha_30_foot:units = "deg" ;
		ted_alpha_30_foot:valid_range = 0., 180. ;
		ted_alpha_30_foot:_Storage = "chunked" ;
		ted_alpha_30_foot:_ChunkSizes = 43200 ;
		ted_alpha_30_foot:_DeflateLevel = 9 ;
		ted_alpha_30_foot:_Shuffle = "true" ;
		ted_alpha_30_foot:_FillValue = -1e+31 ;
	float meped_alpha_0_sat(time) ;
		meped_alpha_0_sat:long_name = "MEPED 0 deg telescope pitch angle (satellite)" ;
		meped_alpha_0_sat:units = "deg" ;
		meped_alpha_0_sat:valid_range = 0., 180. ;
		meped_alpha_0_sat:_Storage = "chunked" ;
		meped_alpha_0_sat:_ChunkSizes = 43200 ;
		meped_alpha_0_sat:_DeflateLevel = 9 ;
		meped_alpha_0_sat:_Shuffle = "true" ;
		meped_alpha_0_sat:_FillValue = -1e+31 ;
	float meped_alpha_90_sat(time) ;
		meped_alpha_90_sat:long_name = "MEPED 90 deg telescope pitch angle (satellite)" ;
		meped_alpha_90_sat:units = "deg" ;
		meped_alpha_90_sat:valid_range = 0., 180. ;
		meped_alpha_90_sat:_Storage = "chunked" ;
		meped_alpha_90_sat:_ChunkSizes = 43200 ;
		meped_alpha_90_sat:_DeflateLevel = 9 ;
		meped_alpha_90_sat:_Shuffle = "true" ;
		meped_alpha_90_sat:_FillValue = -1e+31 ;
	float meped_alpha_0_foot(time) ;
		meped_alpha_0_foot:long_name = "MEPED 0 deg telescope pitch angle (foot of field line)" ;
		meped_alpha_0_foot:units = "deg" ;
		meped_alpha_0_foot:valid_range = 0., 180. ;
		meped_alpha_0_foot:_Storage = "chunked" ;
		meped_alpha_0_foot:_ChunkSizes = 43200 ;
		meped_alpha_0_foot:_DeflateLevel = 9 ;
		meped_alpha_0_foot:_Shuffle = "true" ;
		meped_alpha_0_foot:_FillValue = -1e+31 ;
	float meped_alpha_90_foot(time) ;
		meped_alpha_90_foot:long_name = "MEPED 90 deg telescope pitch angle (foot of field line)" ;
		meped_alpha_90_foot:units = "deg" ;
		meped_alpha_90_foot:valid_range = 0., 180. ;
		meped_alpha_90_foot:_Storage = "chunked" ;
		meped_alpha_90_foot:_ChunkSizes = 43200 ;
		meped_alpha_90_foot:_DeflateLevel = 9 ;
		meped_alpha_90_foot:_Shuffle = "true" ;
		meped_alpha_90_foot:_FillValue = -1e+31 ;
	float L_IGRF(time) ;
		L_IGRF:long_name = "L value from IGRF field" ;
		L_IGRF:units = "" ;
		L_IGRF:valid_range = 0., 20. ;
		L_IGRF:_Storage = "chunked" ;
		L_IGRF:_ChunkSizes = 43200 ;
		L_IGRF:_DeflateLevel = 9 ;
		L_IGRF:_Shuffle = "true" ;
		L_IGRF:_FillValue = -1e+31 ;
	float MLT(time) ;
		MLT:long_name = "Magnetic local time (hours)" ;
		MLT:units = "hours" ;
		MLT:valid_range = 0., 25. ;
		MLT:_Storage = "chunked" ;
		MLT:_ChunkSizes = 43200 ;
		MLT:_DeflateLevel = 9 ;
		MLT:_Shuffle = "true" ;
		MLT:_FillValue = -1e+31 ;
	byte ted_IFC_on(time) ;
		ted_IFC_on:long_name = "TED IFC flag (0 off 1 on)" ;
		ted_IFC_on:units = "on/off" ;
		ted_IFC_on:valid_range = 0., 1. ;
		ted_IFC_on:_Storage = "chunked" ;
		ted_IFC_on:_ChunkSizes = 43200 ;
		ted_IFC_on:_DeflateLevel = 9 ;
		ted_IFC_on:_Shuffle = "true" ;
		ted_IFC_on:_FillValue = -1 ;
	byte mep_IFC_on(time) ;
		mep_IFC_on:long_name = "MEPED IFC flag (0 off 1 on)" ;
		mep_IFC_on:units = "on/off" ;
		mep_IFC_on:valid_range = 0., 1. ;
		mep_IFC_on:_Storage = "chunked" ;
		mep_IFC_on:_ChunkSizes = 43200 ;
		mep_IFC_on:_DeflateLevel = 9 ;
		mep_IFC_on:_Shuffle = "true" ;
		mep_IFC_on:_FillValue = -1 ;

// global attributes:
		:title = "POES/MetOp: Particle Precipitation (These data have known contamination problems. Please consult provider for usage recommendations.)" ;
		:naming_authority = "gov.noaa.ngdc" ;
		:time_coverage_duration = "1day" ;
		:time_coverage_resolution = "2sec" ;
		:geospatial_lat_min = "-90" ;
		:geospatial_lat_max = "90" ;
		:geospatial_lat_unit = "degrees" ;
		:geospatial_lon_min = "0" ;
		:geospatial_lon_max = "360" ;
		:geospatial_lon_units = "degrees East" ;
		:geospatial_vertical_min = "850" ;
		:geospatial_vertical_max = "850" ;
		:geospatial_vertical_units = "km" ;
		:geospatial_vertical_positive = "up" ;
		:point_of_contact = "Rob Redmon" ;
		:institution = "NOAA National Centers for Environmental Information" ;
		:creator = "National Centers for Environmental Information" ;
		:creator_url = "http://www.ngdc.noaa.gov/stp/satellite/poes/index.html" ;
		:creator_email = "Rob.Redmon@noaa.gov" ;
		:publisher_name = "Rob Redmon" ;
		:publisher_url = "http://www.ngdc.noaa.gov/stp/satellite/poes/index.html" ;
		:publisher_email = "Rob.Redmon@noaa.gov" ;
		:release = "Public Release" ;
		:description = "POES/MetOp SEM-2 Data" ;
		:summary = "The POES/MetOp SEM-2 data provide information about the particle radiation surrounding Earth and its effects on the atmosphere" ;
		:keywords_vocabulary = "Earth Science > Sun-earth Interactions > Ionosphere/Magnetosphere Particles > Electron Flux,Earth Science > Sun-earth Interactions > Ionosphere/Magnetosphere Particles " ;
		:comment = "Every effort has been made to provide the highest quality data but the instruments have known inherent limitations. Please contact the data provider for information on how to properly use the data." ;
		:license = "Public" ;
		:Project = "POES/MetOp" ;
		:processing_level = "Level 2, calibrated fluxes" ;
		:_Format = "netCDF-4" ;
}
